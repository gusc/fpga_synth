`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: LU DF (DIP-m)
// Engineer: Tomass Lacis
// 
// Create Date:    19:56:17 06/14/2018 
// Design Name: 
// Module Name:    tableSinewave 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module tableSinewave(idx, sinewave);
parameter USE_UNSIGNED_TABLES = 0;
input [9:0] idx;
output reg [11:0] sinewave = 0;
always @(idx) begin

	if (USE_UNSIGNED_TABLES)
		// Samples: 1024
		// Top value: 4095
		// Mid value: 2047
		// Bottom value: 0
		case(idx)
			0: sinewave = 12'h800; // Dec: 2048
			1: sinewave = 12'h80c; // Dec: 2060
			2: sinewave = 12'h819; // Dec: 2073
			3: sinewave = 12'h825; // Dec: 2085
			4: sinewave = 12'h832; // Dec: 2098
			5: sinewave = 12'h83e; // Dec: 2110
			6: sinewave = 12'h84b; // Dec: 2123
			7: sinewave = 12'h857; // Dec: 2135
			8: sinewave = 12'h864; // Dec: 2148
			9: sinewave = 12'h870; // Dec: 2160
		  10: sinewave = 12'h87d; // Dec: 2173
		  11: sinewave = 12'h88a; // Dec: 2186
		  12: sinewave = 12'h896; // Dec: 2198
		  13: sinewave = 12'h8a3; // Dec: 2211
		  14: sinewave = 12'h8af; // Dec: 2223
		  15: sinewave = 12'h8bc; // Dec: 2236
		  16: sinewave = 12'h8c8; // Dec: 2248
		  17: sinewave = 12'h8d5; // Dec: 2261
		  18: sinewave = 12'h8e1; // Dec: 2273
		  19: sinewave = 12'h8ee; // Dec: 2286
		  20: sinewave = 12'h8fa; // Dec: 2298
		  21: sinewave = 12'h907; // Dec: 2311
		  22: sinewave = 12'h913; // Dec: 2323
		  23: sinewave = 12'h91f; // Dec: 2335
		  24: sinewave = 12'h92c; // Dec: 2348
		  25: sinewave = 12'h938; // Dec: 2360
		  26: sinewave = 12'h945; // Dec: 2373
		  27: sinewave = 12'h951; // Dec: 2385
		  28: sinewave = 12'h95d; // Dec: 2397
		  29: sinewave = 12'h96a; // Dec: 2410
		  30: sinewave = 12'h976; // Dec: 2422
		  31: sinewave = 12'h983; // Dec: 2435
		  32: sinewave = 12'h98f; // Dec: 2447
		  33: sinewave = 12'h99b; // Dec: 2459
		  34: sinewave = 12'h9a7; // Dec: 2471
		  35: sinewave = 12'h9b4; // Dec: 2484
		  36: sinewave = 12'h9c0; // Dec: 2496
		  37: sinewave = 12'h9cc; // Dec: 2508
		  38: sinewave = 12'h9d8; // Dec: 2520
		  39: sinewave = 12'h9e5; // Dec: 2533
		  40: sinewave = 12'h9f1; // Dec: 2545
		  41: sinewave = 12'h9fd; // Dec: 2557
		  42: sinewave = 12'ha09; // Dec: 2569
		  43: sinewave = 12'ha15; // Dec: 2581
		  44: sinewave = 12'ha21; // Dec: 2593
		  45: sinewave = 12'ha2e; // Dec: 2606
		  46: sinewave = 12'ha3a; // Dec: 2618
		  47: sinewave = 12'ha46; // Dec: 2630
		  48: sinewave = 12'ha52; // Dec: 2642
		  49: sinewave = 12'ha5e; // Dec: 2654
		  50: sinewave = 12'ha6a; // Dec: 2666
		  51: sinewave = 12'ha76; // Dec: 2678
		  52: sinewave = 12'ha82; // Dec: 2690
		  53: sinewave = 12'ha8e; // Dec: 2702
		  54: sinewave = 12'ha99; // Dec: 2713
		  55: sinewave = 12'haa5; // Dec: 2725
		  56: sinewave = 12'hab1; // Dec: 2737
		  57: sinewave = 12'habd; // Dec: 2749
		  58: sinewave = 12'hac9; // Dec: 2761
		  59: sinewave = 12'had4; // Dec: 2772
		  60: sinewave = 12'hae0; // Dec: 2784
		  61: sinewave = 12'haec; // Dec: 2796
		  62: sinewave = 12'haf8; // Dec: 2808
		  63: sinewave = 12'hb03; // Dec: 2819
		  64: sinewave = 12'hb0f; // Dec: 2831
		  65: sinewave = 12'hb1a; // Dec: 2842
		  66: sinewave = 12'hb26; // Dec: 2854
		  67: sinewave = 12'hb32; // Dec: 2866
		  68: sinewave = 12'hb3d; // Dec: 2877
		  69: sinewave = 12'hb48; // Dec: 2888
		  70: sinewave = 12'hb54; // Dec: 2900
		  71: sinewave = 12'hb5f; // Dec: 2911
		  72: sinewave = 12'hb6b; // Dec: 2923
		  73: sinewave = 12'hb76; // Dec: 2934
		  74: sinewave = 12'hb81; // Dec: 2945
		  75: sinewave = 12'hb8d; // Dec: 2957
		  76: sinewave = 12'hb98; // Dec: 2968
		  77: sinewave = 12'hba3; // Dec: 2979
		  78: sinewave = 12'hbae; // Dec: 2990
		  79: sinewave = 12'hbb9; // Dec: 3001
		  80: sinewave = 12'hbc4; // Dec: 3012
		  81: sinewave = 12'hbd0; // Dec: 3024
		  82: sinewave = 12'hbdb; // Dec: 3035
		  83: sinewave = 12'hbe6; // Dec: 3046
		  84: sinewave = 12'hbf0; // Dec: 3056
		  85: sinewave = 12'hbfb; // Dec: 3067
		  86: sinewave = 12'hc06; // Dec: 3078
		  87: sinewave = 12'hc11; // Dec: 3089
		  88: sinewave = 12'hc1c; // Dec: 3100
		  89: sinewave = 12'hc27; // Dec: 3111
		  90: sinewave = 12'hc31; // Dec: 3121
		  91: sinewave = 12'hc3c; // Dec: 3132
		  92: sinewave = 12'hc47; // Dec: 3143
		  93: sinewave = 12'hc51; // Dec: 3153
		  94: sinewave = 12'hc5c; // Dec: 3164
		  95: sinewave = 12'hc66; // Dec: 3174
		  96: sinewave = 12'hc71; // Dec: 3185
		  97: sinewave = 12'hc7b; // Dec: 3195
		  98: sinewave = 12'hc86; // Dec: 3206
		  99: sinewave = 12'hc90; // Dec: 3216
		 100: sinewave = 12'hc9a; // Dec: 3226
		 101: sinewave = 12'hca4; // Dec: 3236
		 102: sinewave = 12'hcaf; // Dec: 3247
		 103: sinewave = 12'hcb9; // Dec: 3257
		 104: sinewave = 12'hcc3; // Dec: 3267
		 105: sinewave = 12'hccd; // Dec: 3277
		 106: sinewave = 12'hcd7; // Dec: 3287
		 107: sinewave = 12'hce1; // Dec: 3297
		 108: sinewave = 12'hceb; // Dec: 3307
		 109: sinewave = 12'hcf5; // Dec: 3317
		 110: sinewave = 12'hcff; // Dec: 3327
		 111: sinewave = 12'hd08; // Dec: 3336
		 112: sinewave = 12'hd12; // Dec: 3346
		 113: sinewave = 12'hd1c; // Dec: 3356
		 114: sinewave = 12'hd25; // Dec: 3365
		 115: sinewave = 12'hd2f; // Dec: 3375
		 116: sinewave = 12'hd39; // Dec: 3385
		 117: sinewave = 12'hd42; // Dec: 3394
		 118: sinewave = 12'hd4b; // Dec: 3403
		 119: sinewave = 12'hd55; // Dec: 3413
		 120: sinewave = 12'hd5e; // Dec: 3422
		 121: sinewave = 12'hd67; // Dec: 3431
		 122: sinewave = 12'hd71; // Dec: 3441
		 123: sinewave = 12'hd7a; // Dec: 3450
		 124: sinewave = 12'hd83; // Dec: 3459
		 125: sinewave = 12'hd8c; // Dec: 3468
		 126: sinewave = 12'hd95; // Dec: 3477
		 127: sinewave = 12'hd9e; // Dec: 3486
		 128: sinewave = 12'hda7; // Dec: 3495
		 129: sinewave = 12'hdb0; // Dec: 3504
		 130: sinewave = 12'hdb9; // Dec: 3513
		 131: sinewave = 12'hdc1; // Dec: 3521
		 132: sinewave = 12'hdca; // Dec: 3530
		 133: sinewave = 12'hdd3; // Dec: 3539
		 134: sinewave = 12'hddb; // Dec: 3547
		 135: sinewave = 12'hde4; // Dec: 3556
		 136: sinewave = 12'hdec; // Dec: 3564
		 137: sinewave = 12'hdf5; // Dec: 3573
		 138: sinewave = 12'hdfd; // Dec: 3581
		 139: sinewave = 12'he05; // Dec: 3589
		 140: sinewave = 12'he0e; // Dec: 3598
		 141: sinewave = 12'he16; // Dec: 3606
		 142: sinewave = 12'he1e; // Dec: 3614
		 143: sinewave = 12'he26; // Dec: 3622
		 144: sinewave = 12'he2e; // Dec: 3630
		 145: sinewave = 12'he36; // Dec: 3638
		 146: sinewave = 12'he3e; // Dec: 3646
		 147: sinewave = 12'he45; // Dec: 3653
		 148: sinewave = 12'he4d; // Dec: 3661
		 149: sinewave = 12'he55; // Dec: 3669
		 150: sinewave = 12'he5d; // Dec: 3677
		 151: sinewave = 12'he64; // Dec: 3684
		 152: sinewave = 12'he6c; // Dec: 3692
		 153: sinewave = 12'he73; // Dec: 3699
		 154: sinewave = 12'he7b; // Dec: 3707
		 155: sinewave = 12'he82; // Dec: 3714
		 156: sinewave = 12'he89; // Dec: 3721
		 157: sinewave = 12'he90; // Dec: 3728
		 158: sinewave = 12'he97; // Dec: 3735
		 159: sinewave = 12'he9f; // Dec: 3743
		 160: sinewave = 12'hea6; // Dec: 3750
		 161: sinewave = 12'heac; // Dec: 3756
		 162: sinewave = 12'heb3; // Dec: 3763
		 163: sinewave = 12'heba; // Dec: 3770
		 164: sinewave = 12'hec1; // Dec: 3777
		 165: sinewave = 12'hec8; // Dec: 3784
		 166: sinewave = 12'hece; // Dec: 3790
		 167: sinewave = 12'hed5; // Dec: 3797
		 168: sinewave = 12'hedb; // Dec: 3803
		 169: sinewave = 12'hee2; // Dec: 3810
		 170: sinewave = 12'hee8; // Dec: 3816
		 171: sinewave = 12'heee; // Dec: 3822
		 172: sinewave = 12'hef5; // Dec: 3829
		 173: sinewave = 12'hefb; // Dec: 3835
		 174: sinewave = 12'hf01; // Dec: 3841
		 175: sinewave = 12'hf07; // Dec: 3847
		 176: sinewave = 12'hf0d; // Dec: 3853
		 177: sinewave = 12'hf13; // Dec: 3859
		 178: sinewave = 12'hf18; // Dec: 3864
		 179: sinewave = 12'hf1e; // Dec: 3870
		 180: sinewave = 12'hf24; // Dec: 3876
		 181: sinewave = 12'hf2a; // Dec: 3882
		 182: sinewave = 12'hf2f; // Dec: 3887
		 183: sinewave = 12'hf35; // Dec: 3893
		 184: sinewave = 12'hf3a; // Dec: 3898
		 185: sinewave = 12'hf3f; // Dec: 3903
		 186: sinewave = 12'hf45; // Dec: 3909
		 187: sinewave = 12'hf4a; // Dec: 3914
		 188: sinewave = 12'hf4f; // Dec: 3919
		 189: sinewave = 12'hf54; // Dec: 3924
		 190: sinewave = 12'hf59; // Dec: 3929
		 191: sinewave = 12'hf5e; // Dec: 3934
		 192: sinewave = 12'hf63; // Dec: 3939
		 193: sinewave = 12'hf67; // Dec: 3943
		 194: sinewave = 12'hf6c; // Dec: 3948
		 195: sinewave = 12'hf71; // Dec: 3953
		 196: sinewave = 12'hf75; // Dec: 3957
		 197: sinewave = 12'hf7a; // Dec: 3962
		 198: sinewave = 12'hf7e; // Dec: 3966
		 199: sinewave = 12'hf83; // Dec: 3971
		 200: sinewave = 12'hf87; // Dec: 3975
		 201: sinewave = 12'hf8b; // Dec: 3979
		 202: sinewave = 12'hf8f; // Dec: 3983
		 203: sinewave = 12'hf93; // Dec: 3987
		 204: sinewave = 12'hf97; // Dec: 3991
		 205: sinewave = 12'hf9b; // Dec: 3995
		 206: sinewave = 12'hf9f; // Dec: 3999
		 207: sinewave = 12'hfa3; // Dec: 4003
		 208: sinewave = 12'hfa6; // Dec: 4006
		 209: sinewave = 12'hfaa; // Dec: 4010
		 210: sinewave = 12'hfae; // Dec: 4014
		 211: sinewave = 12'hfb1; // Dec: 4017
		 212: sinewave = 12'hfb4; // Dec: 4020
		 213: sinewave = 12'hfb8; // Dec: 4024
		 214: sinewave = 12'hfbb; // Dec: 4027
		 215: sinewave = 12'hfbe; // Dec: 4030
		 216: sinewave = 12'hfc1; // Dec: 4033
		 217: sinewave = 12'hfc4; // Dec: 4036
		 218: sinewave = 12'hfc7; // Dec: 4039
		 219: sinewave = 12'hfca; // Dec: 4042
		 220: sinewave = 12'hfcd; // Dec: 4045
		 221: sinewave = 12'hfcf; // Dec: 4047
		 222: sinewave = 12'hfd2; // Dec: 4050
		 223: sinewave = 12'hfd5; // Dec: 4053
		 224: sinewave = 12'hfd7; // Dec: 4055
		 225: sinewave = 12'hfda; // Dec: 4058
		 226: sinewave = 12'hfdc; // Dec: 4060
		 227: sinewave = 12'hfde; // Dec: 4062
		 228: sinewave = 12'hfe0; // Dec: 4064
		 229: sinewave = 12'hfe2; // Dec: 4066
		 230: sinewave = 12'hfe5; // Dec: 4069
		 231: sinewave = 12'hfe6; // Dec: 4070
		 232: sinewave = 12'hfe8; // Dec: 4072
		 233: sinewave = 12'hfea; // Dec: 4074
		 234: sinewave = 12'hfec; // Dec: 4076
		 235: sinewave = 12'hfee; // Dec: 4078
		 236: sinewave = 12'hfef; // Dec: 4079
		 237: sinewave = 12'hff1; // Dec: 4081
		 238: sinewave = 12'hff2; // Dec: 4082
		 239: sinewave = 12'hff3; // Dec: 4083
		 240: sinewave = 12'hff5; // Dec: 4085
		 241: sinewave = 12'hff6; // Dec: 4086
		 242: sinewave = 12'hff7; // Dec: 4087
		 243: sinewave = 12'hff8; // Dec: 4088
		 244: sinewave = 12'hff9; // Dec: 4089
		 245: sinewave = 12'hffa; // Dec: 4090
		 246: sinewave = 12'hffb; // Dec: 4091
		 247: sinewave = 12'hffb; // Dec: 4091
		 248: sinewave = 12'hffc; // Dec: 4092
		 249: sinewave = 12'hffd; // Dec: 4093
		 250: sinewave = 12'hffd; // Dec: 4093
		 251: sinewave = 12'hffe; // Dec: 4094
		 252: sinewave = 12'hffe; // Dec: 4094
		 253: sinewave = 12'hffe; // Dec: 4094
		 254: sinewave = 12'hffe; // Dec: 4094
		 255: sinewave = 12'hffe; // Dec: 4094
		 256: sinewave = 12'hfff; // Dec: 4095
		 257: sinewave = 12'hffe; // Dec: 4094
		 258: sinewave = 12'hffe; // Dec: 4094
		 259: sinewave = 12'hffe; // Dec: 4094
		 260: sinewave = 12'hffe; // Dec: 4094
		 261: sinewave = 12'hffe; // Dec: 4094
		 262: sinewave = 12'hffd; // Dec: 4093
		 263: sinewave = 12'hffd; // Dec: 4093
		 264: sinewave = 12'hffc; // Dec: 4092
		 265: sinewave = 12'hffb; // Dec: 4091
		 266: sinewave = 12'hffb; // Dec: 4091
		 267: sinewave = 12'hffa; // Dec: 4090
		 268: sinewave = 12'hff9; // Dec: 4089
		 269: sinewave = 12'hff8; // Dec: 4088
		 270: sinewave = 12'hff7; // Dec: 4087
		 271: sinewave = 12'hff6; // Dec: 4086
		 272: sinewave = 12'hff5; // Dec: 4085
		 273: sinewave = 12'hff3; // Dec: 4083
		 274: sinewave = 12'hff2; // Dec: 4082
		 275: sinewave = 12'hff1; // Dec: 4081
		 276: sinewave = 12'hfef; // Dec: 4079
		 277: sinewave = 12'hfee; // Dec: 4078
		 278: sinewave = 12'hfec; // Dec: 4076
		 279: sinewave = 12'hfea; // Dec: 4074
		 280: sinewave = 12'hfe8; // Dec: 4072
		 281: sinewave = 12'hfe6; // Dec: 4070
		 282: sinewave = 12'hfe5; // Dec: 4069
		 283: sinewave = 12'hfe2; // Dec: 4066
		 284: sinewave = 12'hfe0; // Dec: 4064
		 285: sinewave = 12'hfde; // Dec: 4062
		 286: sinewave = 12'hfdc; // Dec: 4060
		 287: sinewave = 12'hfda; // Dec: 4058
		 288: sinewave = 12'hfd7; // Dec: 4055
		 289: sinewave = 12'hfd5; // Dec: 4053
		 290: sinewave = 12'hfd2; // Dec: 4050
		 291: sinewave = 12'hfcf; // Dec: 4047
		 292: sinewave = 12'hfcd; // Dec: 4045
		 293: sinewave = 12'hfca; // Dec: 4042
		 294: sinewave = 12'hfc7; // Dec: 4039
		 295: sinewave = 12'hfc4; // Dec: 4036
		 296: sinewave = 12'hfc1; // Dec: 4033
		 297: sinewave = 12'hfbe; // Dec: 4030
		 298: sinewave = 12'hfbb; // Dec: 4027
		 299: sinewave = 12'hfb8; // Dec: 4024
		 300: sinewave = 12'hfb4; // Dec: 4020
		 301: sinewave = 12'hfb1; // Dec: 4017
		 302: sinewave = 12'hfae; // Dec: 4014
		 303: sinewave = 12'hfaa; // Dec: 4010
		 304: sinewave = 12'hfa6; // Dec: 4006
		 305: sinewave = 12'hfa3; // Dec: 4003
		 306: sinewave = 12'hf9f; // Dec: 3999
		 307: sinewave = 12'hf9b; // Dec: 3995
		 308: sinewave = 12'hf97; // Dec: 3991
		 309: sinewave = 12'hf93; // Dec: 3987
		 310: sinewave = 12'hf8f; // Dec: 3983
		 311: sinewave = 12'hf8b; // Dec: 3979
		 312: sinewave = 12'hf87; // Dec: 3975
		 313: sinewave = 12'hf83; // Dec: 3971
		 314: sinewave = 12'hf7e; // Dec: 3966
		 315: sinewave = 12'hf7a; // Dec: 3962
		 316: sinewave = 12'hf75; // Dec: 3957
		 317: sinewave = 12'hf71; // Dec: 3953
		 318: sinewave = 12'hf6c; // Dec: 3948
		 319: sinewave = 12'hf67; // Dec: 3943
		 320: sinewave = 12'hf63; // Dec: 3939
		 321: sinewave = 12'hf5e; // Dec: 3934
		 322: sinewave = 12'hf59; // Dec: 3929
		 323: sinewave = 12'hf54; // Dec: 3924
		 324: sinewave = 12'hf4f; // Dec: 3919
		 325: sinewave = 12'hf4a; // Dec: 3914
		 326: sinewave = 12'hf45; // Dec: 3909
		 327: sinewave = 12'hf3f; // Dec: 3903
		 328: sinewave = 12'hf3a; // Dec: 3898
		 329: sinewave = 12'hf35; // Dec: 3893
		 330: sinewave = 12'hf2f; // Dec: 3887
		 331: sinewave = 12'hf2a; // Dec: 3882
		 332: sinewave = 12'hf24; // Dec: 3876
		 333: sinewave = 12'hf1e; // Dec: 3870
		 334: sinewave = 12'hf18; // Dec: 3864
		 335: sinewave = 12'hf13; // Dec: 3859
		 336: sinewave = 12'hf0d; // Dec: 3853
		 337: sinewave = 12'hf07; // Dec: 3847
		 338: sinewave = 12'hf01; // Dec: 3841
		 339: sinewave = 12'hefb; // Dec: 3835
		 340: sinewave = 12'hef5; // Dec: 3829
		 341: sinewave = 12'heee; // Dec: 3822
		 342: sinewave = 12'hee8; // Dec: 3816
		 343: sinewave = 12'hee2; // Dec: 3810
		 344: sinewave = 12'hedb; // Dec: 3803
		 345: sinewave = 12'hed5; // Dec: 3797
		 346: sinewave = 12'hece; // Dec: 3790
		 347: sinewave = 12'hec8; // Dec: 3784
		 348: sinewave = 12'hec1; // Dec: 3777
		 349: sinewave = 12'heba; // Dec: 3770
		 350: sinewave = 12'heb3; // Dec: 3763
		 351: sinewave = 12'heac; // Dec: 3756
		 352: sinewave = 12'hea6; // Dec: 3750
		 353: sinewave = 12'he9f; // Dec: 3743
		 354: sinewave = 12'he97; // Dec: 3735
		 355: sinewave = 12'he90; // Dec: 3728
		 356: sinewave = 12'he89; // Dec: 3721
		 357: sinewave = 12'he82; // Dec: 3714
		 358: sinewave = 12'he7b; // Dec: 3707
		 359: sinewave = 12'he73; // Dec: 3699
		 360: sinewave = 12'he6c; // Dec: 3692
		 361: sinewave = 12'he64; // Dec: 3684
		 362: sinewave = 12'he5d; // Dec: 3677
		 363: sinewave = 12'he55; // Dec: 3669
		 364: sinewave = 12'he4d; // Dec: 3661
		 365: sinewave = 12'he45; // Dec: 3653
		 366: sinewave = 12'he3e; // Dec: 3646
		 367: sinewave = 12'he36; // Dec: 3638
		 368: sinewave = 12'he2e; // Dec: 3630
		 369: sinewave = 12'he26; // Dec: 3622
		 370: sinewave = 12'he1e; // Dec: 3614
		 371: sinewave = 12'he16; // Dec: 3606
		 372: sinewave = 12'he0e; // Dec: 3598
		 373: sinewave = 12'he05; // Dec: 3589
		 374: sinewave = 12'hdfd; // Dec: 3581
		 375: sinewave = 12'hdf5; // Dec: 3573
		 376: sinewave = 12'hdec; // Dec: 3564
		 377: sinewave = 12'hde4; // Dec: 3556
		 378: sinewave = 12'hddb; // Dec: 3547
		 379: sinewave = 12'hdd3; // Dec: 3539
		 380: sinewave = 12'hdca; // Dec: 3530
		 381: sinewave = 12'hdc1; // Dec: 3521
		 382: sinewave = 12'hdb9; // Dec: 3513
		 383: sinewave = 12'hdb0; // Dec: 3504
		 384: sinewave = 12'hda7; // Dec: 3495
		 385: sinewave = 12'hd9e; // Dec: 3486
		 386: sinewave = 12'hd95; // Dec: 3477
		 387: sinewave = 12'hd8c; // Dec: 3468
		 388: sinewave = 12'hd83; // Dec: 3459
		 389: sinewave = 12'hd7a; // Dec: 3450
		 390: sinewave = 12'hd71; // Dec: 3441
		 391: sinewave = 12'hd67; // Dec: 3431
		 392: sinewave = 12'hd5e; // Dec: 3422
		 393: sinewave = 12'hd55; // Dec: 3413
		 394: sinewave = 12'hd4b; // Dec: 3403
		 395: sinewave = 12'hd42; // Dec: 3394
		 396: sinewave = 12'hd39; // Dec: 3385
		 397: sinewave = 12'hd2f; // Dec: 3375
		 398: sinewave = 12'hd25; // Dec: 3365
		 399: sinewave = 12'hd1c; // Dec: 3356
		 400: sinewave = 12'hd12; // Dec: 3346
		 401: sinewave = 12'hd08; // Dec: 3336
		 402: sinewave = 12'hcff; // Dec: 3327
		 403: sinewave = 12'hcf5; // Dec: 3317
		 404: sinewave = 12'hceb; // Dec: 3307
		 405: sinewave = 12'hce1; // Dec: 3297
		 406: sinewave = 12'hcd7; // Dec: 3287
		 407: sinewave = 12'hccd; // Dec: 3277
		 408: sinewave = 12'hcc3; // Dec: 3267
		 409: sinewave = 12'hcb9; // Dec: 3257
		 410: sinewave = 12'hcaf; // Dec: 3247
		 411: sinewave = 12'hca4; // Dec: 3236
		 412: sinewave = 12'hc9a; // Dec: 3226
		 413: sinewave = 12'hc90; // Dec: 3216
		 414: sinewave = 12'hc86; // Dec: 3206
		 415: sinewave = 12'hc7b; // Dec: 3195
		 416: sinewave = 12'hc71; // Dec: 3185
		 417: sinewave = 12'hc66; // Dec: 3174
		 418: sinewave = 12'hc5c; // Dec: 3164
		 419: sinewave = 12'hc51; // Dec: 3153
		 420: sinewave = 12'hc47; // Dec: 3143
		 421: sinewave = 12'hc3c; // Dec: 3132
		 422: sinewave = 12'hc31; // Dec: 3121
		 423: sinewave = 12'hc27; // Dec: 3111
		 424: sinewave = 12'hc1c; // Dec: 3100
		 425: sinewave = 12'hc11; // Dec: 3089
		 426: sinewave = 12'hc06; // Dec: 3078
		 427: sinewave = 12'hbfb; // Dec: 3067
		 428: sinewave = 12'hbf0; // Dec: 3056
		 429: sinewave = 12'hbe6; // Dec: 3046
		 430: sinewave = 12'hbdb; // Dec: 3035
		 431: sinewave = 12'hbd0; // Dec: 3024
		 432: sinewave = 12'hbc4; // Dec: 3012
		 433: sinewave = 12'hbb9; // Dec: 3001
		 434: sinewave = 12'hbae; // Dec: 2990
		 435: sinewave = 12'hba3; // Dec: 2979
		 436: sinewave = 12'hb98; // Dec: 2968
		 437: sinewave = 12'hb8d; // Dec: 2957
		 438: sinewave = 12'hb81; // Dec: 2945
		 439: sinewave = 12'hb76; // Dec: 2934
		 440: sinewave = 12'hb6b; // Dec: 2923
		 441: sinewave = 12'hb5f; // Dec: 2911
		 442: sinewave = 12'hb54; // Dec: 2900
		 443: sinewave = 12'hb48; // Dec: 2888
		 444: sinewave = 12'hb3d; // Dec: 2877
		 445: sinewave = 12'hb32; // Dec: 2866
		 446: sinewave = 12'hb26; // Dec: 2854
		 447: sinewave = 12'hb1a; // Dec: 2842
		 448: sinewave = 12'hb0f; // Dec: 2831
		 449: sinewave = 12'hb03; // Dec: 2819
		 450: sinewave = 12'haf8; // Dec: 2808
		 451: sinewave = 12'haec; // Dec: 2796
		 452: sinewave = 12'hae0; // Dec: 2784
		 453: sinewave = 12'had4; // Dec: 2772
		 454: sinewave = 12'hac9; // Dec: 2761
		 455: sinewave = 12'habd; // Dec: 2749
		 456: sinewave = 12'hab1; // Dec: 2737
		 457: sinewave = 12'haa5; // Dec: 2725
		 458: sinewave = 12'ha99; // Dec: 2713
		 459: sinewave = 12'ha8e; // Dec: 2702
		 460: sinewave = 12'ha82; // Dec: 2690
		 461: sinewave = 12'ha76; // Dec: 2678
		 462: sinewave = 12'ha6a; // Dec: 2666
		 463: sinewave = 12'ha5e; // Dec: 2654
		 464: sinewave = 12'ha52; // Dec: 2642
		 465: sinewave = 12'ha46; // Dec: 2630
		 466: sinewave = 12'ha3a; // Dec: 2618
		 467: sinewave = 12'ha2e; // Dec: 2606
		 468: sinewave = 12'ha21; // Dec: 2593
		 469: sinewave = 12'ha15; // Dec: 2581
		 470: sinewave = 12'ha09; // Dec: 2569
		 471: sinewave = 12'h9fd; // Dec: 2557
		 472: sinewave = 12'h9f1; // Dec: 2545
		 473: sinewave = 12'h9e5; // Dec: 2533
		 474: sinewave = 12'h9d8; // Dec: 2520
		 475: sinewave = 12'h9cc; // Dec: 2508
		 476: sinewave = 12'h9c0; // Dec: 2496
		 477: sinewave = 12'h9b4; // Dec: 2484
		 478: sinewave = 12'h9a7; // Dec: 2471
		 479: sinewave = 12'h99b; // Dec: 2459
		 480: sinewave = 12'h98f; // Dec: 2447
		 481: sinewave = 12'h983; // Dec: 2435
		 482: sinewave = 12'h976; // Dec: 2422
		 483: sinewave = 12'h96a; // Dec: 2410
		 484: sinewave = 12'h95d; // Dec: 2397
		 485: sinewave = 12'h951; // Dec: 2385
		 486: sinewave = 12'h945; // Dec: 2373
		 487: sinewave = 12'h938; // Dec: 2360
		 488: sinewave = 12'h92c; // Dec: 2348
		 489: sinewave = 12'h91f; // Dec: 2335
		 490: sinewave = 12'h913; // Dec: 2323
		 491: sinewave = 12'h907; // Dec: 2311
		 492: sinewave = 12'h8fa; // Dec: 2298
		 493: sinewave = 12'h8ee; // Dec: 2286
		 494: sinewave = 12'h8e1; // Dec: 2273
		 495: sinewave = 12'h8d5; // Dec: 2261
		 496: sinewave = 12'h8c8; // Dec: 2248
		 497: sinewave = 12'h8bc; // Dec: 2236
		 498: sinewave = 12'h8af; // Dec: 2223
		 499: sinewave = 12'h8a3; // Dec: 2211
		 500: sinewave = 12'h896; // Dec: 2198
		 501: sinewave = 12'h88a; // Dec: 2186
		 502: sinewave = 12'h87d; // Dec: 2173
		 503: sinewave = 12'h870; // Dec: 2160
		 504: sinewave = 12'h864; // Dec: 2148
		 505: sinewave = 12'h857; // Dec: 2135
		 506: sinewave = 12'h84b; // Dec: 2123
		 507: sinewave = 12'h83e; // Dec: 2110
		 508: sinewave = 12'h832; // Dec: 2098
		 509: sinewave = 12'h825; // Dec: 2085
		 510: sinewave = 12'h819; // Dec: 2073
		 511: sinewave = 12'h80c; // Dec: 2060
		 512: sinewave = 12'h800; // Dec: 2048
		 513: sinewave = 12'h7f3; // Dec: 2035
		 514: sinewave = 12'h7e6; // Dec: 2022
		 515: sinewave = 12'h7da; // Dec: 2010
		 516: sinewave = 12'h7cd; // Dec: 1997
		 517: sinewave = 12'h7c1; // Dec: 1985
		 518: sinewave = 12'h7b4; // Dec: 1972
		 519: sinewave = 12'h7a8; // Dec: 1960
		 520: sinewave = 12'h79b; // Dec: 1947
		 521: sinewave = 12'h78f; // Dec: 1935
		 522: sinewave = 12'h782; // Dec: 1922
		 523: sinewave = 12'h775; // Dec: 1909
		 524: sinewave = 12'h769; // Dec: 1897
		 525: sinewave = 12'h75c; // Dec: 1884
		 526: sinewave = 12'h750; // Dec: 1872
		 527: sinewave = 12'h743; // Dec: 1859
		 528: sinewave = 12'h737; // Dec: 1847
		 529: sinewave = 12'h72a; // Dec: 1834
		 530: sinewave = 12'h71e; // Dec: 1822
		 531: sinewave = 12'h711; // Dec: 1809
		 532: sinewave = 12'h705; // Dec: 1797
		 533: sinewave = 12'h6f8; // Dec: 1784
		 534: sinewave = 12'h6ec; // Dec: 1772
		 535: sinewave = 12'h6e0; // Dec: 1760
		 536: sinewave = 12'h6d3; // Dec: 1747
		 537: sinewave = 12'h6c7; // Dec: 1735
		 538: sinewave = 12'h6ba; // Dec: 1722
		 539: sinewave = 12'h6ae; // Dec: 1710
		 540: sinewave = 12'h6a2; // Dec: 1698
		 541: sinewave = 12'h695; // Dec: 1685
		 542: sinewave = 12'h689; // Dec: 1673
		 543: sinewave = 12'h67c; // Dec: 1660
		 544: sinewave = 12'h670; // Dec: 1648
		 545: sinewave = 12'h664; // Dec: 1636
		 546: sinewave = 12'h658; // Dec: 1624
		 547: sinewave = 12'h64b; // Dec: 1611
		 548: sinewave = 12'h63f; // Dec: 1599
		 549: sinewave = 12'h633; // Dec: 1587
		 550: sinewave = 12'h627; // Dec: 1575
		 551: sinewave = 12'h61a; // Dec: 1562
		 552: sinewave = 12'h60e; // Dec: 1550
		 553: sinewave = 12'h602; // Dec: 1538
		 554: sinewave = 12'h5f6; // Dec: 1526
		 555: sinewave = 12'h5ea; // Dec: 1514
		 556: sinewave = 12'h5de; // Dec: 1502
		 557: sinewave = 12'h5d1; // Dec: 1489
		 558: sinewave = 12'h5c5; // Dec: 1477
		 559: sinewave = 12'h5b9; // Dec: 1465
		 560: sinewave = 12'h5ad; // Dec: 1453
		 561: sinewave = 12'h5a1; // Dec: 1441
		 562: sinewave = 12'h595; // Dec: 1429
		 563: sinewave = 12'h589; // Dec: 1417
		 564: sinewave = 12'h57d; // Dec: 1405
		 565: sinewave = 12'h571; // Dec: 1393
		 566: sinewave = 12'h566; // Dec: 1382
		 567: sinewave = 12'h55a; // Dec: 1370
		 568: sinewave = 12'h54e; // Dec: 1358
		 569: sinewave = 12'h542; // Dec: 1346
		 570: sinewave = 12'h536; // Dec: 1334
		 571: sinewave = 12'h52b; // Dec: 1323
		 572: sinewave = 12'h51f; // Dec: 1311
		 573: sinewave = 12'h513; // Dec: 1299
		 574: sinewave = 12'h507; // Dec: 1287
		 575: sinewave = 12'h4fc; // Dec: 1276
		 576: sinewave = 12'h4f0; // Dec: 1264
		 577: sinewave = 12'h4e5; // Dec: 1253
		 578: sinewave = 12'h4d9; // Dec: 1241
		 579: sinewave = 12'h4cd; // Dec: 1229
		 580: sinewave = 12'h4c2; // Dec: 1218
		 581: sinewave = 12'h4b7; // Dec: 1207
		 582: sinewave = 12'h4ab; // Dec: 1195
		 583: sinewave = 12'h4a0; // Dec: 1184
		 584: sinewave = 12'h494; // Dec: 1172
		 585: sinewave = 12'h489; // Dec: 1161
		 586: sinewave = 12'h47e; // Dec: 1150
		 587: sinewave = 12'h472; // Dec: 1138
		 588: sinewave = 12'h467; // Dec: 1127
		 589: sinewave = 12'h45c; // Dec: 1116
		 590: sinewave = 12'h451; // Dec: 1105
		 591: sinewave = 12'h446; // Dec: 1094
		 592: sinewave = 12'h43b; // Dec: 1083
		 593: sinewave = 12'h42f; // Dec: 1071
		 594: sinewave = 12'h424; // Dec: 1060
		 595: sinewave = 12'h419; // Dec: 1049
		 596: sinewave = 12'h40f; // Dec: 1039
		 597: sinewave = 12'h404; // Dec: 1028
		 598: sinewave = 12'h3f9; // Dec: 1017
		 599: sinewave = 12'h3ee; // Dec: 1006
		 600: sinewave = 12'h3e3; // Dec: 995
		 601: sinewave = 12'h3d8; // Dec: 984
		 602: sinewave = 12'h3ce; // Dec: 974
		 603: sinewave = 12'h3c3; // Dec: 963
		 604: sinewave = 12'h3b8; // Dec: 952
		 605: sinewave = 12'h3ae; // Dec: 942
		 606: sinewave = 12'h3a3; // Dec: 931
		 607: sinewave = 12'h399; // Dec: 921
		 608: sinewave = 12'h38e; // Dec: 910
		 609: sinewave = 12'h384; // Dec: 900
		 610: sinewave = 12'h379; // Dec: 889
		 611: sinewave = 12'h36f; // Dec: 879
		 612: sinewave = 12'h365; // Dec: 869
		 613: sinewave = 12'h35b; // Dec: 859
		 614: sinewave = 12'h350; // Dec: 848
		 615: sinewave = 12'h346; // Dec: 838
		 616: sinewave = 12'h33c; // Dec: 828
		 617: sinewave = 12'h332; // Dec: 818
		 618: sinewave = 12'h328; // Dec: 808
		 619: sinewave = 12'h31e; // Dec: 798
		 620: sinewave = 12'h314; // Dec: 788
		 621: sinewave = 12'h30a; // Dec: 778
		 622: sinewave = 12'h300; // Dec: 768
		 623: sinewave = 12'h2f7; // Dec: 759
		 624: sinewave = 12'h2ed; // Dec: 749
		 625: sinewave = 12'h2e3; // Dec: 739
		 626: sinewave = 12'h2da; // Dec: 730
		 627: sinewave = 12'h2d0; // Dec: 720
		 628: sinewave = 12'h2c6; // Dec: 710
		 629: sinewave = 12'h2bd; // Dec: 701
		 630: sinewave = 12'h2b4; // Dec: 692
		 631: sinewave = 12'h2aa; // Dec: 682
		 632: sinewave = 12'h2a1; // Dec: 673
		 633: sinewave = 12'h298; // Dec: 664
		 634: sinewave = 12'h28e; // Dec: 654
		 635: sinewave = 12'h285; // Dec: 645
		 636: sinewave = 12'h27c; // Dec: 636
		 637: sinewave = 12'h273; // Dec: 627
		 638: sinewave = 12'h26a; // Dec: 618
		 639: sinewave = 12'h261; // Dec: 609
		 640: sinewave = 12'h258; // Dec: 600
		 641: sinewave = 12'h24f; // Dec: 591
		 642: sinewave = 12'h246; // Dec: 582
		 643: sinewave = 12'h23e; // Dec: 574
		 644: sinewave = 12'h235; // Dec: 565
		 645: sinewave = 12'h22c; // Dec: 556
		 646: sinewave = 12'h224; // Dec: 548
		 647: sinewave = 12'h21b; // Dec: 539
		 648: sinewave = 12'h213; // Dec: 531
		 649: sinewave = 12'h20a; // Dec: 522
		 650: sinewave = 12'h202; // Dec: 514
		 651: sinewave = 12'h1fa; // Dec: 506
		 652: sinewave = 12'h1f1; // Dec: 497
		 653: sinewave = 12'h1e9; // Dec: 489
		 654: sinewave = 12'h1e1; // Dec: 481
		 655: sinewave = 12'h1d9; // Dec: 473
		 656: sinewave = 12'h1d1; // Dec: 465
		 657: sinewave = 12'h1c9; // Dec: 457
		 658: sinewave = 12'h1c1; // Dec: 449
		 659: sinewave = 12'h1ba; // Dec: 442
		 660: sinewave = 12'h1b2; // Dec: 434
		 661: sinewave = 12'h1aa; // Dec: 426
		 662: sinewave = 12'h1a2; // Dec: 418
		 663: sinewave = 12'h19b; // Dec: 411
		 664: sinewave = 12'h193; // Dec: 403
		 665: sinewave = 12'h18c; // Dec: 396
		 666: sinewave = 12'h184; // Dec: 388
		 667: sinewave = 12'h17d; // Dec: 381
		 668: sinewave = 12'h176; // Dec: 374
		 669: sinewave = 12'h16f; // Dec: 367
		 670: sinewave = 12'h168; // Dec: 360
		 671: sinewave = 12'h160; // Dec: 352
		 672: sinewave = 12'h159; // Dec: 345
		 673: sinewave = 12'h153; // Dec: 339
		 674: sinewave = 12'h14c; // Dec: 332
		 675: sinewave = 12'h145; // Dec: 325
		 676: sinewave = 12'h13e; // Dec: 318
		 677: sinewave = 12'h137; // Dec: 311
		 678: sinewave = 12'h131; // Dec: 305
		 679: sinewave = 12'h12a; // Dec: 298
		 680: sinewave = 12'h124; // Dec: 292
		 681: sinewave = 12'h11d; // Dec: 285
		 682: sinewave = 12'h117; // Dec: 279
		 683: sinewave = 12'h111; // Dec: 273
		 684: sinewave = 12'h10a; // Dec: 266
		 685: sinewave = 12'h104; // Dec: 260
		 686: sinewave = 12'hfe; // Dec: 254
		 687: sinewave = 12'hf8; // Dec: 248
		 688: sinewave = 12'hf2; // Dec: 242
		 689: sinewave = 12'hec; // Dec: 236
		 690: sinewave = 12'he7; // Dec: 231
		 691: sinewave = 12'he1; // Dec: 225
		 692: sinewave = 12'hdb; // Dec: 219
		 693: sinewave = 12'hd5; // Dec: 213
		 694: sinewave = 12'hd0; // Dec: 208
		 695: sinewave = 12'hca; // Dec: 202
		 696: sinewave = 12'hc5; // Dec: 197
		 697: sinewave = 12'hc0; // Dec: 192
		 698: sinewave = 12'hba; // Dec: 186
		 699: sinewave = 12'hb5; // Dec: 181
		 700: sinewave = 12'hb0; // Dec: 176
		 701: sinewave = 12'hab; // Dec: 171
		 702: sinewave = 12'ha6; // Dec: 166
		 703: sinewave = 12'ha1; // Dec: 161
		 704: sinewave = 12'h9c; // Dec: 156
		 705: sinewave = 12'h98; // Dec: 152
		 706: sinewave = 12'h93; // Dec: 147
		 707: sinewave = 12'h8e; // Dec: 142
		 708: sinewave = 12'h8a; // Dec: 138
		 709: sinewave = 12'h85; // Dec: 133
		 710: sinewave = 12'h81; // Dec: 129
		 711: sinewave = 12'h7c; // Dec: 124
		 712: sinewave = 12'h78; // Dec: 120
		 713: sinewave = 12'h74; // Dec: 116
		 714: sinewave = 12'h70; // Dec: 112
		 715: sinewave = 12'h6c; // Dec: 108
		 716: sinewave = 12'h68; // Dec: 104
		 717: sinewave = 12'h64; // Dec: 100
		 718: sinewave = 12'h60; // Dec: 96
		 719: sinewave = 12'h5c; // Dec: 92
		 720: sinewave = 12'h59; // Dec: 89
		 721: sinewave = 12'h55; // Dec: 85
		 722: sinewave = 12'h51; // Dec: 81
		 723: sinewave = 12'h4e; // Dec: 78
		 724: sinewave = 12'h4b; // Dec: 75
		 725: sinewave = 12'h47; // Dec: 71
		 726: sinewave = 12'h44; // Dec: 68
		 727: sinewave = 12'h41; // Dec: 65
		 728: sinewave = 12'h3e; // Dec: 62
		 729: sinewave = 12'h3b; // Dec: 59
		 730: sinewave = 12'h38; // Dec: 56
		 731: sinewave = 12'h35; // Dec: 53
		 732: sinewave = 12'h32; // Dec: 50
		 733: sinewave = 12'h30; // Dec: 48
		 734: sinewave = 12'h2d; // Dec: 45
		 735: sinewave = 12'h2a; // Dec: 42
		 736: sinewave = 12'h28; // Dec: 40
		 737: sinewave = 12'h25; // Dec: 37
		 738: sinewave = 12'h23; // Dec: 35
		 739: sinewave = 12'h21; // Dec: 33
		 740: sinewave = 12'h1f; // Dec: 31
		 741: sinewave = 12'h1d; // Dec: 29
		 742: sinewave = 12'h1a; // Dec: 26
		 743: sinewave = 12'h19; // Dec: 25
		 744: sinewave = 12'h17; // Dec: 23
		 745: sinewave = 12'h15; // Dec: 21
		 746: sinewave = 12'h13; // Dec: 19
		 747: sinewave = 12'h11; // Dec: 17
		 748: sinewave = 12'h10; // Dec: 16
		 749: sinewave = 12'h0e; // Dec: 14
		 750: sinewave = 12'h0d; // Dec: 13
		 751: sinewave = 12'h0c; // Dec: 12
		 752: sinewave = 12'h0a; // Dec: 10
		 753: sinewave = 12'h09; // Dec: 9
		 754: sinewave = 12'h08; // Dec: 8
		 755: sinewave = 12'h07; // Dec: 7
		 756: sinewave = 12'h06; // Dec: 6
		 757: sinewave = 12'h05; // Dec: 5
		 758: sinewave = 12'h04; // Dec: 4
		 759: sinewave = 12'h04; // Dec: 4
		 760: sinewave = 12'h03; // Dec: 3
		 761: sinewave = 12'h02; // Dec: 2
		 762: sinewave = 12'h02; // Dec: 2
		 763: sinewave = 12'h01; // Dec: 1
		 764: sinewave = 12'h01; // Dec: 1
		 765: sinewave = 12'h01; // Dec: 1
		 766: sinewave = 12'h01; // Dec: 1
		 767: sinewave = 12'h01; // Dec: 1
		 768: sinewave = 12'h00; // Dec: 0
		 769: sinewave = 12'h01; // Dec: 1
		 770: sinewave = 12'h01; // Dec: 1
		 771: sinewave = 12'h01; // Dec: 1
		 772: sinewave = 12'h01; // Dec: 1
		 773: sinewave = 12'h01; // Dec: 1
		 774: sinewave = 12'h02; // Dec: 2
		 775: sinewave = 12'h02; // Dec: 2
		 776: sinewave = 12'h03; // Dec: 3
		 777: sinewave = 12'h04; // Dec: 4
		 778: sinewave = 12'h04; // Dec: 4
		 779: sinewave = 12'h05; // Dec: 5
		 780: sinewave = 12'h06; // Dec: 6
		 781: sinewave = 12'h07; // Dec: 7
		 782: sinewave = 12'h08; // Dec: 8
		 783: sinewave = 12'h09; // Dec: 9
		 784: sinewave = 12'h0a; // Dec: 10
		 785: sinewave = 12'h0c; // Dec: 12
		 786: sinewave = 12'h0d; // Dec: 13
		 787: sinewave = 12'h0e; // Dec: 14
		 788: sinewave = 12'h10; // Dec: 16
		 789: sinewave = 12'h11; // Dec: 17
		 790: sinewave = 12'h13; // Dec: 19
		 791: sinewave = 12'h15; // Dec: 21
		 792: sinewave = 12'h17; // Dec: 23
		 793: sinewave = 12'h19; // Dec: 25
		 794: sinewave = 12'h1a; // Dec: 26
		 795: sinewave = 12'h1d; // Dec: 29
		 796: sinewave = 12'h1f; // Dec: 31
		 797: sinewave = 12'h21; // Dec: 33
		 798: sinewave = 12'h23; // Dec: 35
		 799: sinewave = 12'h25; // Dec: 37
		 800: sinewave = 12'h28; // Dec: 40
		 801: sinewave = 12'h2a; // Dec: 42
		 802: sinewave = 12'h2d; // Dec: 45
		 803: sinewave = 12'h30; // Dec: 48
		 804: sinewave = 12'h32; // Dec: 50
		 805: sinewave = 12'h35; // Dec: 53
		 806: sinewave = 12'h38; // Dec: 56
		 807: sinewave = 12'h3b; // Dec: 59
		 808: sinewave = 12'h3e; // Dec: 62
		 809: sinewave = 12'h41; // Dec: 65
		 810: sinewave = 12'h44; // Dec: 68
		 811: sinewave = 12'h47; // Dec: 71
		 812: sinewave = 12'h4b; // Dec: 75
		 813: sinewave = 12'h4e; // Dec: 78
		 814: sinewave = 12'h51; // Dec: 81
		 815: sinewave = 12'h55; // Dec: 85
		 816: sinewave = 12'h59; // Dec: 89
		 817: sinewave = 12'h5c; // Dec: 92
		 818: sinewave = 12'h60; // Dec: 96
		 819: sinewave = 12'h64; // Dec: 100
		 820: sinewave = 12'h68; // Dec: 104
		 821: sinewave = 12'h6c; // Dec: 108
		 822: sinewave = 12'h70; // Dec: 112
		 823: sinewave = 12'h74; // Dec: 116
		 824: sinewave = 12'h78; // Dec: 120
		 825: sinewave = 12'h7c; // Dec: 124
		 826: sinewave = 12'h81; // Dec: 129
		 827: sinewave = 12'h85; // Dec: 133
		 828: sinewave = 12'h8a; // Dec: 138
		 829: sinewave = 12'h8e; // Dec: 142
		 830: sinewave = 12'h93; // Dec: 147
		 831: sinewave = 12'h98; // Dec: 152
		 832: sinewave = 12'h9c; // Dec: 156
		 833: sinewave = 12'ha1; // Dec: 161
		 834: sinewave = 12'ha6; // Dec: 166
		 835: sinewave = 12'hab; // Dec: 171
		 836: sinewave = 12'hb0; // Dec: 176
		 837: sinewave = 12'hb5; // Dec: 181
		 838: sinewave = 12'hba; // Dec: 186
		 839: sinewave = 12'hc0; // Dec: 192
		 840: sinewave = 12'hc5; // Dec: 197
		 841: sinewave = 12'hca; // Dec: 202
		 842: sinewave = 12'hd0; // Dec: 208
		 843: sinewave = 12'hd5; // Dec: 213
		 844: sinewave = 12'hdb; // Dec: 219
		 845: sinewave = 12'he1; // Dec: 225
		 846: sinewave = 12'he7; // Dec: 231
		 847: sinewave = 12'hec; // Dec: 236
		 848: sinewave = 12'hf2; // Dec: 242
		 849: sinewave = 12'hf8; // Dec: 248
		 850: sinewave = 12'hfe; // Dec: 254
		 851: sinewave = 12'h104; // Dec: 260
		 852: sinewave = 12'h10a; // Dec: 266
		 853: sinewave = 12'h111; // Dec: 273
		 854: sinewave = 12'h117; // Dec: 279
		 855: sinewave = 12'h11d; // Dec: 285
		 856: sinewave = 12'h124; // Dec: 292
		 857: sinewave = 12'h12a; // Dec: 298
		 858: sinewave = 12'h131; // Dec: 305
		 859: sinewave = 12'h137; // Dec: 311
		 860: sinewave = 12'h13e; // Dec: 318
		 861: sinewave = 12'h145; // Dec: 325
		 862: sinewave = 12'h14c; // Dec: 332
		 863: sinewave = 12'h153; // Dec: 339
		 864: sinewave = 12'h159; // Dec: 345
		 865: sinewave = 12'h160; // Dec: 352
		 866: sinewave = 12'h168; // Dec: 360
		 867: sinewave = 12'h16f; // Dec: 367
		 868: sinewave = 12'h176; // Dec: 374
		 869: sinewave = 12'h17d; // Dec: 381
		 870: sinewave = 12'h184; // Dec: 388
		 871: sinewave = 12'h18c; // Dec: 396
		 872: sinewave = 12'h193; // Dec: 403
		 873: sinewave = 12'h19b; // Dec: 411
		 874: sinewave = 12'h1a2; // Dec: 418
		 875: sinewave = 12'h1aa; // Dec: 426
		 876: sinewave = 12'h1b2; // Dec: 434
		 877: sinewave = 12'h1ba; // Dec: 442
		 878: sinewave = 12'h1c1; // Dec: 449
		 879: sinewave = 12'h1c9; // Dec: 457
		 880: sinewave = 12'h1d1; // Dec: 465
		 881: sinewave = 12'h1d9; // Dec: 473
		 882: sinewave = 12'h1e1; // Dec: 481
		 883: sinewave = 12'h1e9; // Dec: 489
		 884: sinewave = 12'h1f1; // Dec: 497
		 885: sinewave = 12'h1fa; // Dec: 506
		 886: sinewave = 12'h202; // Dec: 514
		 887: sinewave = 12'h20a; // Dec: 522
		 888: sinewave = 12'h213; // Dec: 531
		 889: sinewave = 12'h21b; // Dec: 539
		 890: sinewave = 12'h224; // Dec: 548
		 891: sinewave = 12'h22c; // Dec: 556
		 892: sinewave = 12'h235; // Dec: 565
		 893: sinewave = 12'h23e; // Dec: 574
		 894: sinewave = 12'h246; // Dec: 582
		 895: sinewave = 12'h24f; // Dec: 591
		 896: sinewave = 12'h258; // Dec: 600
		 897: sinewave = 12'h261; // Dec: 609
		 898: sinewave = 12'h26a; // Dec: 618
		 899: sinewave = 12'h273; // Dec: 627
		 900: sinewave = 12'h27c; // Dec: 636
		 901: sinewave = 12'h285; // Dec: 645
		 902: sinewave = 12'h28e; // Dec: 654
		 903: sinewave = 12'h298; // Dec: 664
		 904: sinewave = 12'h2a1; // Dec: 673
		 905: sinewave = 12'h2aa; // Dec: 682
		 906: sinewave = 12'h2b4; // Dec: 692
		 907: sinewave = 12'h2bd; // Dec: 701
		 908: sinewave = 12'h2c6; // Dec: 710
		 909: sinewave = 12'h2d0; // Dec: 720
		 910: sinewave = 12'h2da; // Dec: 730
		 911: sinewave = 12'h2e3; // Dec: 739
		 912: sinewave = 12'h2ed; // Dec: 749
		 913: sinewave = 12'h2f7; // Dec: 759
		 914: sinewave = 12'h300; // Dec: 768
		 915: sinewave = 12'h30a; // Dec: 778
		 916: sinewave = 12'h314; // Dec: 788
		 917: sinewave = 12'h31e; // Dec: 798
		 918: sinewave = 12'h328; // Dec: 808
		 919: sinewave = 12'h332; // Dec: 818
		 920: sinewave = 12'h33c; // Dec: 828
		 921: sinewave = 12'h346; // Dec: 838
		 922: sinewave = 12'h350; // Dec: 848
		 923: sinewave = 12'h35b; // Dec: 859
		 924: sinewave = 12'h365; // Dec: 869
		 925: sinewave = 12'h36f; // Dec: 879
		 926: sinewave = 12'h379; // Dec: 889
		 927: sinewave = 12'h384; // Dec: 900
		 928: sinewave = 12'h38e; // Dec: 910
		 929: sinewave = 12'h399; // Dec: 921
		 930: sinewave = 12'h3a3; // Dec: 931
		 931: sinewave = 12'h3ae; // Dec: 942
		 932: sinewave = 12'h3b8; // Dec: 952
		 933: sinewave = 12'h3c3; // Dec: 963
		 934: sinewave = 12'h3ce; // Dec: 974
		 935: sinewave = 12'h3d8; // Dec: 984
		 936: sinewave = 12'h3e3; // Dec: 995
		 937: sinewave = 12'h3ee; // Dec: 1006
		 938: sinewave = 12'h3f9; // Dec: 1017
		 939: sinewave = 12'h404; // Dec: 1028
		 940: sinewave = 12'h40f; // Dec: 1039
		 941: sinewave = 12'h419; // Dec: 1049
		 942: sinewave = 12'h424; // Dec: 1060
		 943: sinewave = 12'h42f; // Dec: 1071
		 944: sinewave = 12'h43b; // Dec: 1083
		 945: sinewave = 12'h446; // Dec: 1094
		 946: sinewave = 12'h451; // Dec: 1105
		 947: sinewave = 12'h45c; // Dec: 1116
		 948: sinewave = 12'h467; // Dec: 1127
		 949: sinewave = 12'h472; // Dec: 1138
		 950: sinewave = 12'h47e; // Dec: 1150
		 951: sinewave = 12'h489; // Dec: 1161
		 952: sinewave = 12'h494; // Dec: 1172
		 953: sinewave = 12'h4a0; // Dec: 1184
		 954: sinewave = 12'h4ab; // Dec: 1195
		 955: sinewave = 12'h4b7; // Dec: 1207
		 956: sinewave = 12'h4c2; // Dec: 1218
		 957: sinewave = 12'h4cd; // Dec: 1229
		 958: sinewave = 12'h4d9; // Dec: 1241
		 959: sinewave = 12'h4e5; // Dec: 1253
		 960: sinewave = 12'h4f0; // Dec: 1264
		 961: sinewave = 12'h4fc; // Dec: 1276
		 962: sinewave = 12'h507; // Dec: 1287
		 963: sinewave = 12'h513; // Dec: 1299
		 964: sinewave = 12'h51f; // Dec: 1311
		 965: sinewave = 12'h52b; // Dec: 1323
		 966: sinewave = 12'h536; // Dec: 1334
		 967: sinewave = 12'h542; // Dec: 1346
		 968: sinewave = 12'h54e; // Dec: 1358
		 969: sinewave = 12'h55a; // Dec: 1370
		 970: sinewave = 12'h566; // Dec: 1382
		 971: sinewave = 12'h571; // Dec: 1393
		 972: sinewave = 12'h57d; // Dec: 1405
		 973: sinewave = 12'h589; // Dec: 1417
		 974: sinewave = 12'h595; // Dec: 1429
		 975: sinewave = 12'h5a1; // Dec: 1441
		 976: sinewave = 12'h5ad; // Dec: 1453
		 977: sinewave = 12'h5b9; // Dec: 1465
		 978: sinewave = 12'h5c5; // Dec: 1477
		 979: sinewave = 12'h5d1; // Dec: 1489
		 980: sinewave = 12'h5de; // Dec: 1502
		 981: sinewave = 12'h5ea; // Dec: 1514
		 982: sinewave = 12'h5f6; // Dec: 1526
		 983: sinewave = 12'h602; // Dec: 1538
		 984: sinewave = 12'h60e; // Dec: 1550
		 985: sinewave = 12'h61a; // Dec: 1562
		 986: sinewave = 12'h627; // Dec: 1575
		 987: sinewave = 12'h633; // Dec: 1587
		 988: sinewave = 12'h63f; // Dec: 1599
		 989: sinewave = 12'h64b; // Dec: 1611
		 990: sinewave = 12'h658; // Dec: 1624
		 991: sinewave = 12'h664; // Dec: 1636
		 992: sinewave = 12'h670; // Dec: 1648
		 993: sinewave = 12'h67c; // Dec: 1660
		 994: sinewave = 12'h689; // Dec: 1673
		 995: sinewave = 12'h695; // Dec: 1685
		 996: sinewave = 12'h6a2; // Dec: 1698
		 997: sinewave = 12'h6ae; // Dec: 1710
		 998: sinewave = 12'h6ba; // Dec: 1722
		 999: sinewave = 12'h6c7; // Dec: 1735
		1000: sinewave = 12'h6d3; // Dec: 1747
		1001: sinewave = 12'h6e0; // Dec: 1760
		1002: sinewave = 12'h6ec; // Dec: 1772
		1003: sinewave = 12'h6f8; // Dec: 1784
		1004: sinewave = 12'h705; // Dec: 1797
		1005: sinewave = 12'h711; // Dec: 1809
		1006: sinewave = 12'h71e; // Dec: 1822
		1007: sinewave = 12'h72a; // Dec: 1834
		1008: sinewave = 12'h737; // Dec: 1847
		1009: sinewave = 12'h743; // Dec: 1859
		1010: sinewave = 12'h750; // Dec: 1872
		1011: sinewave = 12'h75c; // Dec: 1884
		1012: sinewave = 12'h769; // Dec: 1897
		1013: sinewave = 12'h775; // Dec: 1909
		1014: sinewave = 12'h782; // Dec: 1922
		1015: sinewave = 12'h78f; // Dec: 1935
		1016: sinewave = 12'h79b; // Dec: 1947
		1017: sinewave = 12'h7a8; // Dec: 1960
		1018: sinewave = 12'h7b4; // Dec: 1972
		1019: sinewave = 12'h7c1; // Dec: 1985
		1020: sinewave = 12'h7cd; // Dec: 1997
		1021: sinewave = 12'h7da; // Dec: 2010
		1022: sinewave = 12'h7e6; // Dec: 2022
		1023: sinewave = 12'h7f3; // Dec: 2035
		endcase		
	else
		// Samples: 1024
		// Top value: 2047
		// Mid value: 0
		// Bottom value: -2047
		case(idx)
			0: sinewave = 12'h00; // Dec: 0
			1: sinewave = 12'h0c; // Dec: 12
			2: sinewave = 12'h19; // Dec: 25
			3: sinewave = 12'h25; // Dec: 37
			4: sinewave = 12'h32; // Dec: 50
			5: sinewave = 12'h3e; // Dec: 62
			6: sinewave = 12'h4b; // Dec: 75
			7: sinewave = 12'h57; // Dec: 87
			8: sinewave = 12'h64; // Dec: 100
			9: sinewave = 12'h70; // Dec: 112
		  10: sinewave = 12'h7d; // Dec: 125
		  11: sinewave = 12'h8a; // Dec: 138
		  12: sinewave = 12'h96; // Dec: 150
		  13: sinewave = 12'ha3; // Dec: 163
		  14: sinewave = 12'haf; // Dec: 175
		  15: sinewave = 12'hbc; // Dec: 188
		  16: sinewave = 12'hc8; // Dec: 200
		  17: sinewave = 12'hd5; // Dec: 213
		  18: sinewave = 12'he1; // Dec: 225
		  19: sinewave = 12'hee; // Dec: 238
		  20: sinewave = 12'hfa; // Dec: 250
		  21: sinewave = 12'h107; // Dec: 263
		  22: sinewave = 12'h113; // Dec: 275
		  23: sinewave = 12'h11f; // Dec: 287
		  24: sinewave = 12'h12c; // Dec: 300
		  25: sinewave = 12'h138; // Dec: 312
		  26: sinewave = 12'h145; // Dec: 325
		  27: sinewave = 12'h151; // Dec: 337
		  28: sinewave = 12'h15d; // Dec: 349
		  29: sinewave = 12'h16a; // Dec: 362
		  30: sinewave = 12'h176; // Dec: 374
		  31: sinewave = 12'h183; // Dec: 387
		  32: sinewave = 12'h18f; // Dec: 399
		  33: sinewave = 12'h19b; // Dec: 411
		  34: sinewave = 12'h1a7; // Dec: 423
		  35: sinewave = 12'h1b4; // Dec: 436
		  36: sinewave = 12'h1c0; // Dec: 448
		  37: sinewave = 12'h1cc; // Dec: 460
		  38: sinewave = 12'h1d8; // Dec: 472
		  39: sinewave = 12'h1e5; // Dec: 485
		  40: sinewave = 12'h1f1; // Dec: 497
		  41: sinewave = 12'h1fd; // Dec: 509
		  42: sinewave = 12'h209; // Dec: 521
		  43: sinewave = 12'h215; // Dec: 533
		  44: sinewave = 12'h221; // Dec: 545
		  45: sinewave = 12'h22e; // Dec: 558
		  46: sinewave = 12'h23a; // Dec: 570
		  47: sinewave = 12'h246; // Dec: 582
		  48: sinewave = 12'h252; // Dec: 594
		  49: sinewave = 12'h25e; // Dec: 606
		  50: sinewave = 12'h26a; // Dec: 618
		  51: sinewave = 12'h276; // Dec: 630
		  52: sinewave = 12'h282; // Dec: 642
		  53: sinewave = 12'h28e; // Dec: 654
		  54: sinewave = 12'h299; // Dec: 665
		  55: sinewave = 12'h2a5; // Dec: 677
		  56: sinewave = 12'h2b1; // Dec: 689
		  57: sinewave = 12'h2bd; // Dec: 701
		  58: sinewave = 12'h2c9; // Dec: 713
		  59: sinewave = 12'h2d4; // Dec: 724
		  60: sinewave = 12'h2e0; // Dec: 736
		  61: sinewave = 12'h2ec; // Dec: 748
		  62: sinewave = 12'h2f8; // Dec: 760
		  63: sinewave = 12'h303; // Dec: 771
		  64: sinewave = 12'h30f; // Dec: 783
		  65: sinewave = 12'h31a; // Dec: 794
		  66: sinewave = 12'h326; // Dec: 806
		  67: sinewave = 12'h332; // Dec: 818
		  68: sinewave = 12'h33d; // Dec: 829
		  69: sinewave = 12'h348; // Dec: 840
		  70: sinewave = 12'h354; // Dec: 852
		  71: sinewave = 12'h35f; // Dec: 863
		  72: sinewave = 12'h36b; // Dec: 875
		  73: sinewave = 12'h376; // Dec: 886
		  74: sinewave = 12'h381; // Dec: 897
		  75: sinewave = 12'h38d; // Dec: 909
		  76: sinewave = 12'h398; // Dec: 920
		  77: sinewave = 12'h3a3; // Dec: 931
		  78: sinewave = 12'h3ae; // Dec: 942
		  79: sinewave = 12'h3b9; // Dec: 953
		  80: sinewave = 12'h3c4; // Dec: 964
		  81: sinewave = 12'h3d0; // Dec: 976
		  82: sinewave = 12'h3db; // Dec: 987
		  83: sinewave = 12'h3e6; // Dec: 998
		  84: sinewave = 12'h3f0; // Dec: 1008
		  85: sinewave = 12'h3fb; // Dec: 1019
		  86: sinewave = 12'h406; // Dec: 1030
		  87: sinewave = 12'h411; // Dec: 1041
		  88: sinewave = 12'h41c; // Dec: 1052
		  89: sinewave = 12'h427; // Dec: 1063
		  90: sinewave = 12'h431; // Dec: 1073
		  91: sinewave = 12'h43c; // Dec: 1084
		  92: sinewave = 12'h447; // Dec: 1095
		  93: sinewave = 12'h451; // Dec: 1105
		  94: sinewave = 12'h45c; // Dec: 1116
		  95: sinewave = 12'h466; // Dec: 1126
		  96: sinewave = 12'h471; // Dec: 1137
		  97: sinewave = 12'h47b; // Dec: 1147
		  98: sinewave = 12'h486; // Dec: 1158
		  99: sinewave = 12'h490; // Dec: 1168
		 100: sinewave = 12'h49a; // Dec: 1178
		 101: sinewave = 12'h4a4; // Dec: 1188
		 102: sinewave = 12'h4af; // Dec: 1199
		 103: sinewave = 12'h4b9; // Dec: 1209
		 104: sinewave = 12'h4c3; // Dec: 1219
		 105: sinewave = 12'h4cd; // Dec: 1229
		 106: sinewave = 12'h4d7; // Dec: 1239
		 107: sinewave = 12'h4e1; // Dec: 1249
		 108: sinewave = 12'h4eb; // Dec: 1259
		 109: sinewave = 12'h4f5; // Dec: 1269
		 110: sinewave = 12'h4ff; // Dec: 1279
		 111: sinewave = 12'h508; // Dec: 1288
		 112: sinewave = 12'h512; // Dec: 1298
		 113: sinewave = 12'h51c; // Dec: 1308
		 114: sinewave = 12'h525; // Dec: 1317
		 115: sinewave = 12'h52f; // Dec: 1327
		 116: sinewave = 12'h539; // Dec: 1337
		 117: sinewave = 12'h542; // Dec: 1346
		 118: sinewave = 12'h54b; // Dec: 1355
		 119: sinewave = 12'h555; // Dec: 1365
		 120: sinewave = 12'h55e; // Dec: 1374
		 121: sinewave = 12'h567; // Dec: 1383
		 122: sinewave = 12'h571; // Dec: 1393
		 123: sinewave = 12'h57a; // Dec: 1402
		 124: sinewave = 12'h583; // Dec: 1411
		 125: sinewave = 12'h58c; // Dec: 1420
		 126: sinewave = 12'h595; // Dec: 1429
		 127: sinewave = 12'h59e; // Dec: 1438
		 128: sinewave = 12'h5a7; // Dec: 1447
		 129: sinewave = 12'h5b0; // Dec: 1456
		 130: sinewave = 12'h5b9; // Dec: 1465
		 131: sinewave = 12'h5c1; // Dec: 1473
		 132: sinewave = 12'h5ca; // Dec: 1482
		 133: sinewave = 12'h5d3; // Dec: 1491
		 134: sinewave = 12'h5db; // Dec: 1499
		 135: sinewave = 12'h5e4; // Dec: 1508
		 136: sinewave = 12'h5ec; // Dec: 1516
		 137: sinewave = 12'h5f5; // Dec: 1525
		 138: sinewave = 12'h5fd; // Dec: 1533
		 139: sinewave = 12'h605; // Dec: 1541
		 140: sinewave = 12'h60e; // Dec: 1550
		 141: sinewave = 12'h616; // Dec: 1558
		 142: sinewave = 12'h61e; // Dec: 1566
		 143: sinewave = 12'h626; // Dec: 1574
		 144: sinewave = 12'h62e; // Dec: 1582
		 145: sinewave = 12'h636; // Dec: 1590
		 146: sinewave = 12'h63e; // Dec: 1598
		 147: sinewave = 12'h645; // Dec: 1605
		 148: sinewave = 12'h64d; // Dec: 1613
		 149: sinewave = 12'h655; // Dec: 1621
		 150: sinewave = 12'h65d; // Dec: 1629
		 151: sinewave = 12'h664; // Dec: 1636
		 152: sinewave = 12'h66c; // Dec: 1644
		 153: sinewave = 12'h673; // Dec: 1651
		 154: sinewave = 12'h67b; // Dec: 1659
		 155: sinewave = 12'h682; // Dec: 1666
		 156: sinewave = 12'h689; // Dec: 1673
		 157: sinewave = 12'h690; // Dec: 1680
		 158: sinewave = 12'h697; // Dec: 1687
		 159: sinewave = 12'h69f; // Dec: 1695
		 160: sinewave = 12'h6a6; // Dec: 1702
		 161: sinewave = 12'h6ac; // Dec: 1708
		 162: sinewave = 12'h6b3; // Dec: 1715
		 163: sinewave = 12'h6ba; // Dec: 1722
		 164: sinewave = 12'h6c1; // Dec: 1729
		 165: sinewave = 12'h6c8; // Dec: 1736
		 166: sinewave = 12'h6ce; // Dec: 1742
		 167: sinewave = 12'h6d5; // Dec: 1749
		 168: sinewave = 12'h6db; // Dec: 1755
		 169: sinewave = 12'h6e2; // Dec: 1762
		 170: sinewave = 12'h6e8; // Dec: 1768
		 171: sinewave = 12'h6ee; // Dec: 1774
		 172: sinewave = 12'h6f5; // Dec: 1781
		 173: sinewave = 12'h6fb; // Dec: 1787
		 174: sinewave = 12'h701; // Dec: 1793
		 175: sinewave = 12'h707; // Dec: 1799
		 176: sinewave = 12'h70d; // Dec: 1805
		 177: sinewave = 12'h713; // Dec: 1811
		 178: sinewave = 12'h718; // Dec: 1816
		 179: sinewave = 12'h71e; // Dec: 1822
		 180: sinewave = 12'h724; // Dec: 1828
		 181: sinewave = 12'h72a; // Dec: 1834
		 182: sinewave = 12'h72f; // Dec: 1839
		 183: sinewave = 12'h735; // Dec: 1845
		 184: sinewave = 12'h73a; // Dec: 1850
		 185: sinewave = 12'h73f; // Dec: 1855
		 186: sinewave = 12'h745; // Dec: 1861
		 187: sinewave = 12'h74a; // Dec: 1866
		 188: sinewave = 12'h74f; // Dec: 1871
		 189: sinewave = 12'h754; // Dec: 1876
		 190: sinewave = 12'h759; // Dec: 1881
		 191: sinewave = 12'h75e; // Dec: 1886
		 192: sinewave = 12'h763; // Dec: 1891
		 193: sinewave = 12'h767; // Dec: 1895
		 194: sinewave = 12'h76c; // Dec: 1900
		 195: sinewave = 12'h771; // Dec: 1905
		 196: sinewave = 12'h775; // Dec: 1909
		 197: sinewave = 12'h77a; // Dec: 1914
		 198: sinewave = 12'h77e; // Dec: 1918
		 199: sinewave = 12'h783; // Dec: 1923
		 200: sinewave = 12'h787; // Dec: 1927
		 201: sinewave = 12'h78b; // Dec: 1931
		 202: sinewave = 12'h78f; // Dec: 1935
		 203: sinewave = 12'h793; // Dec: 1939
		 204: sinewave = 12'h797; // Dec: 1943
		 205: sinewave = 12'h79b; // Dec: 1947
		 206: sinewave = 12'h79f; // Dec: 1951
		 207: sinewave = 12'h7a3; // Dec: 1955
		 208: sinewave = 12'h7a6; // Dec: 1958
		 209: sinewave = 12'h7aa; // Dec: 1962
		 210: sinewave = 12'h7ae; // Dec: 1966
		 211: sinewave = 12'h7b1; // Dec: 1969
		 212: sinewave = 12'h7b4; // Dec: 1972
		 213: sinewave = 12'h7b8; // Dec: 1976
		 214: sinewave = 12'h7bb; // Dec: 1979
		 215: sinewave = 12'h7be; // Dec: 1982
		 216: sinewave = 12'h7c1; // Dec: 1985
		 217: sinewave = 12'h7c4; // Dec: 1988
		 218: sinewave = 12'h7c7; // Dec: 1991
		 219: sinewave = 12'h7ca; // Dec: 1994
		 220: sinewave = 12'h7cd; // Dec: 1997
		 221: sinewave = 12'h7cf; // Dec: 1999
		 222: sinewave = 12'h7d2; // Dec: 2002
		 223: sinewave = 12'h7d5; // Dec: 2005
		 224: sinewave = 12'h7d7; // Dec: 2007
		 225: sinewave = 12'h7da; // Dec: 2010
		 226: sinewave = 12'h7dc; // Dec: 2012
		 227: sinewave = 12'h7de; // Dec: 2014
		 228: sinewave = 12'h7e0; // Dec: 2016
		 229: sinewave = 12'h7e2; // Dec: 2018
		 230: sinewave = 12'h7e5; // Dec: 2021
		 231: sinewave = 12'h7e6; // Dec: 2022
		 232: sinewave = 12'h7e8; // Dec: 2024
		 233: sinewave = 12'h7ea; // Dec: 2026
		 234: sinewave = 12'h7ec; // Dec: 2028
		 235: sinewave = 12'h7ee; // Dec: 2030
		 236: sinewave = 12'h7ef; // Dec: 2031
		 237: sinewave = 12'h7f1; // Dec: 2033
		 238: sinewave = 12'h7f2; // Dec: 2034
		 239: sinewave = 12'h7f3; // Dec: 2035
		 240: sinewave = 12'h7f5; // Dec: 2037
		 241: sinewave = 12'h7f6; // Dec: 2038
		 242: sinewave = 12'h7f7; // Dec: 2039
		 243: sinewave = 12'h7f8; // Dec: 2040
		 244: sinewave = 12'h7f9; // Dec: 2041
		 245: sinewave = 12'h7fa; // Dec: 2042
		 246: sinewave = 12'h7fb; // Dec: 2043
		 247: sinewave = 12'h7fb; // Dec: 2043
		 248: sinewave = 12'h7fc; // Dec: 2044
		 249: sinewave = 12'h7fd; // Dec: 2045
		 250: sinewave = 12'h7fd; // Dec: 2045
		 251: sinewave = 12'h7fe; // Dec: 2046
		 252: sinewave = 12'h7fe; // Dec: 2046
		 253: sinewave = 12'h7fe; // Dec: 2046
		 254: sinewave = 12'h7fe; // Dec: 2046
		 255: sinewave = 12'h7fe; // Dec: 2046
		 256: sinewave = 12'h7ff; // Dec: 2047
		 257: sinewave = 12'h7fe; // Dec: 2046
		 258: sinewave = 12'h7fe; // Dec: 2046
		 259: sinewave = 12'h7fe; // Dec: 2046
		 260: sinewave = 12'h7fe; // Dec: 2046
		 261: sinewave = 12'h7fe; // Dec: 2046
		 262: sinewave = 12'h7fd; // Dec: 2045
		 263: sinewave = 12'h7fd; // Dec: 2045
		 264: sinewave = 12'h7fc; // Dec: 2044
		 265: sinewave = 12'h7fb; // Dec: 2043
		 266: sinewave = 12'h7fb; // Dec: 2043
		 267: sinewave = 12'h7fa; // Dec: 2042
		 268: sinewave = 12'h7f9; // Dec: 2041
		 269: sinewave = 12'h7f8; // Dec: 2040
		 270: sinewave = 12'h7f7; // Dec: 2039
		 271: sinewave = 12'h7f6; // Dec: 2038
		 272: sinewave = 12'h7f5; // Dec: 2037
		 273: sinewave = 12'h7f3; // Dec: 2035
		 274: sinewave = 12'h7f2; // Dec: 2034
		 275: sinewave = 12'h7f1; // Dec: 2033
		 276: sinewave = 12'h7ef; // Dec: 2031
		 277: sinewave = 12'h7ee; // Dec: 2030
		 278: sinewave = 12'h7ec; // Dec: 2028
		 279: sinewave = 12'h7ea; // Dec: 2026
		 280: sinewave = 12'h7e8; // Dec: 2024
		 281: sinewave = 12'h7e6; // Dec: 2022
		 282: sinewave = 12'h7e5; // Dec: 2021
		 283: sinewave = 12'h7e2; // Dec: 2018
		 284: sinewave = 12'h7e0; // Dec: 2016
		 285: sinewave = 12'h7de; // Dec: 2014
		 286: sinewave = 12'h7dc; // Dec: 2012
		 287: sinewave = 12'h7da; // Dec: 2010
		 288: sinewave = 12'h7d7; // Dec: 2007
		 289: sinewave = 12'h7d5; // Dec: 2005
		 290: sinewave = 12'h7d2; // Dec: 2002
		 291: sinewave = 12'h7cf; // Dec: 1999
		 292: sinewave = 12'h7cd; // Dec: 1997
		 293: sinewave = 12'h7ca; // Dec: 1994
		 294: sinewave = 12'h7c7; // Dec: 1991
		 295: sinewave = 12'h7c4; // Dec: 1988
		 296: sinewave = 12'h7c1; // Dec: 1985
		 297: sinewave = 12'h7be; // Dec: 1982
		 298: sinewave = 12'h7bb; // Dec: 1979
		 299: sinewave = 12'h7b8; // Dec: 1976
		 300: sinewave = 12'h7b4; // Dec: 1972
		 301: sinewave = 12'h7b1; // Dec: 1969
		 302: sinewave = 12'h7ae; // Dec: 1966
		 303: sinewave = 12'h7aa; // Dec: 1962
		 304: sinewave = 12'h7a6; // Dec: 1958
		 305: sinewave = 12'h7a3; // Dec: 1955
		 306: sinewave = 12'h79f; // Dec: 1951
		 307: sinewave = 12'h79b; // Dec: 1947
		 308: sinewave = 12'h797; // Dec: 1943
		 309: sinewave = 12'h793; // Dec: 1939
		 310: sinewave = 12'h78f; // Dec: 1935
		 311: sinewave = 12'h78b; // Dec: 1931
		 312: sinewave = 12'h787; // Dec: 1927
		 313: sinewave = 12'h783; // Dec: 1923
		 314: sinewave = 12'h77e; // Dec: 1918
		 315: sinewave = 12'h77a; // Dec: 1914
		 316: sinewave = 12'h775; // Dec: 1909
		 317: sinewave = 12'h771; // Dec: 1905
		 318: sinewave = 12'h76c; // Dec: 1900
		 319: sinewave = 12'h767; // Dec: 1895
		 320: sinewave = 12'h763; // Dec: 1891
		 321: sinewave = 12'h75e; // Dec: 1886
		 322: sinewave = 12'h759; // Dec: 1881
		 323: sinewave = 12'h754; // Dec: 1876
		 324: sinewave = 12'h74f; // Dec: 1871
		 325: sinewave = 12'h74a; // Dec: 1866
		 326: sinewave = 12'h745; // Dec: 1861
		 327: sinewave = 12'h73f; // Dec: 1855
		 328: sinewave = 12'h73a; // Dec: 1850
		 329: sinewave = 12'h735; // Dec: 1845
		 330: sinewave = 12'h72f; // Dec: 1839
		 331: sinewave = 12'h72a; // Dec: 1834
		 332: sinewave = 12'h724; // Dec: 1828
		 333: sinewave = 12'h71e; // Dec: 1822
		 334: sinewave = 12'h718; // Dec: 1816
		 335: sinewave = 12'h713; // Dec: 1811
		 336: sinewave = 12'h70d; // Dec: 1805
		 337: sinewave = 12'h707; // Dec: 1799
		 338: sinewave = 12'h701; // Dec: 1793
		 339: sinewave = 12'h6fb; // Dec: 1787
		 340: sinewave = 12'h6f5; // Dec: 1781
		 341: sinewave = 12'h6ee; // Dec: 1774
		 342: sinewave = 12'h6e8; // Dec: 1768
		 343: sinewave = 12'h6e2; // Dec: 1762
		 344: sinewave = 12'h6db; // Dec: 1755
		 345: sinewave = 12'h6d5; // Dec: 1749
		 346: sinewave = 12'h6ce; // Dec: 1742
		 347: sinewave = 12'h6c8; // Dec: 1736
		 348: sinewave = 12'h6c1; // Dec: 1729
		 349: sinewave = 12'h6ba; // Dec: 1722
		 350: sinewave = 12'h6b3; // Dec: 1715
		 351: sinewave = 12'h6ac; // Dec: 1708
		 352: sinewave = 12'h6a6; // Dec: 1702
		 353: sinewave = 12'h69f; // Dec: 1695
		 354: sinewave = 12'h697; // Dec: 1687
		 355: sinewave = 12'h690; // Dec: 1680
		 356: sinewave = 12'h689; // Dec: 1673
		 357: sinewave = 12'h682; // Dec: 1666
		 358: sinewave = 12'h67b; // Dec: 1659
		 359: sinewave = 12'h673; // Dec: 1651
		 360: sinewave = 12'h66c; // Dec: 1644
		 361: sinewave = 12'h664; // Dec: 1636
		 362: sinewave = 12'h65d; // Dec: 1629
		 363: sinewave = 12'h655; // Dec: 1621
		 364: sinewave = 12'h64d; // Dec: 1613
		 365: sinewave = 12'h645; // Dec: 1605
		 366: sinewave = 12'h63e; // Dec: 1598
		 367: sinewave = 12'h636; // Dec: 1590
		 368: sinewave = 12'h62e; // Dec: 1582
		 369: sinewave = 12'h626; // Dec: 1574
		 370: sinewave = 12'h61e; // Dec: 1566
		 371: sinewave = 12'h616; // Dec: 1558
		 372: sinewave = 12'h60e; // Dec: 1550
		 373: sinewave = 12'h605; // Dec: 1541
		 374: sinewave = 12'h5fd; // Dec: 1533
		 375: sinewave = 12'h5f5; // Dec: 1525
		 376: sinewave = 12'h5ec; // Dec: 1516
		 377: sinewave = 12'h5e4; // Dec: 1508
		 378: sinewave = 12'h5db; // Dec: 1499
		 379: sinewave = 12'h5d3; // Dec: 1491
		 380: sinewave = 12'h5ca; // Dec: 1482
		 381: sinewave = 12'h5c1; // Dec: 1473
		 382: sinewave = 12'h5b9; // Dec: 1465
		 383: sinewave = 12'h5b0; // Dec: 1456
		 384: sinewave = 12'h5a7; // Dec: 1447
		 385: sinewave = 12'h59e; // Dec: 1438
		 386: sinewave = 12'h595; // Dec: 1429
		 387: sinewave = 12'h58c; // Dec: 1420
		 388: sinewave = 12'h583; // Dec: 1411
		 389: sinewave = 12'h57a; // Dec: 1402
		 390: sinewave = 12'h571; // Dec: 1393
		 391: sinewave = 12'h567; // Dec: 1383
		 392: sinewave = 12'h55e; // Dec: 1374
		 393: sinewave = 12'h555; // Dec: 1365
		 394: sinewave = 12'h54b; // Dec: 1355
		 395: sinewave = 12'h542; // Dec: 1346
		 396: sinewave = 12'h539; // Dec: 1337
		 397: sinewave = 12'h52f; // Dec: 1327
		 398: sinewave = 12'h525; // Dec: 1317
		 399: sinewave = 12'h51c; // Dec: 1308
		 400: sinewave = 12'h512; // Dec: 1298
		 401: sinewave = 12'h508; // Dec: 1288
		 402: sinewave = 12'h4ff; // Dec: 1279
		 403: sinewave = 12'h4f5; // Dec: 1269
		 404: sinewave = 12'h4eb; // Dec: 1259
		 405: sinewave = 12'h4e1; // Dec: 1249
		 406: sinewave = 12'h4d7; // Dec: 1239
		 407: sinewave = 12'h4cd; // Dec: 1229
		 408: sinewave = 12'h4c3; // Dec: 1219
		 409: sinewave = 12'h4b9; // Dec: 1209
		 410: sinewave = 12'h4af; // Dec: 1199
		 411: sinewave = 12'h4a4; // Dec: 1188
		 412: sinewave = 12'h49a; // Dec: 1178
		 413: sinewave = 12'h490; // Dec: 1168
		 414: sinewave = 12'h486; // Dec: 1158
		 415: sinewave = 12'h47b; // Dec: 1147
		 416: sinewave = 12'h471; // Dec: 1137
		 417: sinewave = 12'h466; // Dec: 1126
		 418: sinewave = 12'h45c; // Dec: 1116
		 419: sinewave = 12'h451; // Dec: 1105
		 420: sinewave = 12'h447; // Dec: 1095
		 421: sinewave = 12'h43c; // Dec: 1084
		 422: sinewave = 12'h431; // Dec: 1073
		 423: sinewave = 12'h427; // Dec: 1063
		 424: sinewave = 12'h41c; // Dec: 1052
		 425: sinewave = 12'h411; // Dec: 1041
		 426: sinewave = 12'h406; // Dec: 1030
		 427: sinewave = 12'h3fb; // Dec: 1019
		 428: sinewave = 12'h3f0; // Dec: 1008
		 429: sinewave = 12'h3e6; // Dec: 998
		 430: sinewave = 12'h3db; // Dec: 987
		 431: sinewave = 12'h3d0; // Dec: 976
		 432: sinewave = 12'h3c4; // Dec: 964
		 433: sinewave = 12'h3b9; // Dec: 953
		 434: sinewave = 12'h3ae; // Dec: 942
		 435: sinewave = 12'h3a3; // Dec: 931
		 436: sinewave = 12'h398; // Dec: 920
		 437: sinewave = 12'h38d; // Dec: 909
		 438: sinewave = 12'h381; // Dec: 897
		 439: sinewave = 12'h376; // Dec: 886
		 440: sinewave = 12'h36b; // Dec: 875
		 441: sinewave = 12'h35f; // Dec: 863
		 442: sinewave = 12'h354; // Dec: 852
		 443: sinewave = 12'h348; // Dec: 840
		 444: sinewave = 12'h33d; // Dec: 829
		 445: sinewave = 12'h332; // Dec: 818
		 446: sinewave = 12'h326; // Dec: 806
		 447: sinewave = 12'h31a; // Dec: 794
		 448: sinewave = 12'h30f; // Dec: 783
		 449: sinewave = 12'h303; // Dec: 771
		 450: sinewave = 12'h2f8; // Dec: 760
		 451: sinewave = 12'h2ec; // Dec: 748
		 452: sinewave = 12'h2e0; // Dec: 736
		 453: sinewave = 12'h2d4; // Dec: 724
		 454: sinewave = 12'h2c9; // Dec: 713
		 455: sinewave = 12'h2bd; // Dec: 701
		 456: sinewave = 12'h2b1; // Dec: 689
		 457: sinewave = 12'h2a5; // Dec: 677
		 458: sinewave = 12'h299; // Dec: 665
		 459: sinewave = 12'h28e; // Dec: 654
		 460: sinewave = 12'h282; // Dec: 642
		 461: sinewave = 12'h276; // Dec: 630
		 462: sinewave = 12'h26a; // Dec: 618
		 463: sinewave = 12'h25e; // Dec: 606
		 464: sinewave = 12'h252; // Dec: 594
		 465: sinewave = 12'h246; // Dec: 582
		 466: sinewave = 12'h23a; // Dec: 570
		 467: sinewave = 12'h22e; // Dec: 558
		 468: sinewave = 12'h221; // Dec: 545
		 469: sinewave = 12'h215; // Dec: 533
		 470: sinewave = 12'h209; // Dec: 521
		 471: sinewave = 12'h1fd; // Dec: 509
		 472: sinewave = 12'h1f1; // Dec: 497
		 473: sinewave = 12'h1e5; // Dec: 485
		 474: sinewave = 12'h1d8; // Dec: 472
		 475: sinewave = 12'h1cc; // Dec: 460
		 476: sinewave = 12'h1c0; // Dec: 448
		 477: sinewave = 12'h1b4; // Dec: 436
		 478: sinewave = 12'h1a7; // Dec: 423
		 479: sinewave = 12'h19b; // Dec: 411
		 480: sinewave = 12'h18f; // Dec: 399
		 481: sinewave = 12'h183; // Dec: 387
		 482: sinewave = 12'h176; // Dec: 374
		 483: sinewave = 12'h16a; // Dec: 362
		 484: sinewave = 12'h15d; // Dec: 349
		 485: sinewave = 12'h151; // Dec: 337
		 486: sinewave = 12'h145; // Dec: 325
		 487: sinewave = 12'h138; // Dec: 312
		 488: sinewave = 12'h12c; // Dec: 300
		 489: sinewave = 12'h11f; // Dec: 287
		 490: sinewave = 12'h113; // Dec: 275
		 491: sinewave = 12'h107; // Dec: 263
		 492: sinewave = 12'hfa; // Dec: 250
		 493: sinewave = 12'hee; // Dec: 238
		 494: sinewave = 12'he1; // Dec: 225
		 495: sinewave = 12'hd5; // Dec: 213
		 496: sinewave = 12'hc8; // Dec: 200
		 497: sinewave = 12'hbc; // Dec: 188
		 498: sinewave = 12'haf; // Dec: 175
		 499: sinewave = 12'ha3; // Dec: 163
		 500: sinewave = 12'h96; // Dec: 150
		 501: sinewave = 12'h8a; // Dec: 138
		 502: sinewave = 12'h7d; // Dec: 125
		 503: sinewave = 12'h70; // Dec: 112
		 504: sinewave = 12'h64; // Dec: 100
		 505: sinewave = 12'h57; // Dec: 87
		 506: sinewave = 12'h4b; // Dec: 75
		 507: sinewave = 12'h3e; // Dec: 62
		 508: sinewave = 12'h32; // Dec: 50
		 509: sinewave = 12'h25; // Dec: 37
		 510: sinewave = 12'h19; // Dec: 25
		 511: sinewave = 12'h0c; // Dec: 12
		 512: sinewave = 12'h00; // Dec: 0
		 513: sinewave = 12'hff4; // Dec: -12
		 514: sinewave = 12'hfe7; // Dec: -25
		 515: sinewave = 12'hfdb; // Dec: -37
		 516: sinewave = 12'hfce; // Dec: -50
		 517: sinewave = 12'hfc2; // Dec: -62
		 518: sinewave = 12'hfb5; // Dec: -75
		 519: sinewave = 12'hfa9; // Dec: -87
		 520: sinewave = 12'hf9c; // Dec: -100
		 521: sinewave = 12'hf90; // Dec: -112
		 522: sinewave = 12'hf83; // Dec: -125
		 523: sinewave = 12'hf76; // Dec: -138
		 524: sinewave = 12'hf6a; // Dec: -150
		 525: sinewave = 12'hf5d; // Dec: -163
		 526: sinewave = 12'hf51; // Dec: -175
		 527: sinewave = 12'hf44; // Dec: -188
		 528: sinewave = 12'hf38; // Dec: -200
		 529: sinewave = 12'hf2b; // Dec: -213
		 530: sinewave = 12'hf1f; // Dec: -225
		 531: sinewave = 12'hf12; // Dec: -238
		 532: sinewave = 12'hf06; // Dec: -250
		 533: sinewave = 12'hef9; // Dec: -263
		 534: sinewave = 12'heed; // Dec: -275
		 535: sinewave = 12'hee1; // Dec: -287
		 536: sinewave = 12'hed4; // Dec: -300
		 537: sinewave = 12'hec8; // Dec: -312
		 538: sinewave = 12'hebb; // Dec: -325
		 539: sinewave = 12'heaf; // Dec: -337
		 540: sinewave = 12'hea3; // Dec: -349
		 541: sinewave = 12'he96; // Dec: -362
		 542: sinewave = 12'he8a; // Dec: -374
		 543: sinewave = 12'he7d; // Dec: -387
		 544: sinewave = 12'he71; // Dec: -399
		 545: sinewave = 12'he65; // Dec: -411
		 546: sinewave = 12'he59; // Dec: -423
		 547: sinewave = 12'he4c; // Dec: -436
		 548: sinewave = 12'he40; // Dec: -448
		 549: sinewave = 12'he34; // Dec: -460
		 550: sinewave = 12'he28; // Dec: -472
		 551: sinewave = 12'he1b; // Dec: -485
		 552: sinewave = 12'he0f; // Dec: -497
		 553: sinewave = 12'he03; // Dec: -509
		 554: sinewave = 12'hdf7; // Dec: -521
		 555: sinewave = 12'hdeb; // Dec: -533
		 556: sinewave = 12'hddf; // Dec: -545
		 557: sinewave = 12'hdd2; // Dec: -558
		 558: sinewave = 12'hdc6; // Dec: -570
		 559: sinewave = 12'hdba; // Dec: -582
		 560: sinewave = 12'hdae; // Dec: -594
		 561: sinewave = 12'hda2; // Dec: -606
		 562: sinewave = 12'hd96; // Dec: -618
		 563: sinewave = 12'hd8a; // Dec: -630
		 564: sinewave = 12'hd7e; // Dec: -642
		 565: sinewave = 12'hd72; // Dec: -654
		 566: sinewave = 12'hd67; // Dec: -665
		 567: sinewave = 12'hd5b; // Dec: -677
		 568: sinewave = 12'hd4f; // Dec: -689
		 569: sinewave = 12'hd43; // Dec: -701
		 570: sinewave = 12'hd37; // Dec: -713
		 571: sinewave = 12'hd2c; // Dec: -724
		 572: sinewave = 12'hd20; // Dec: -736
		 573: sinewave = 12'hd14; // Dec: -748
		 574: sinewave = 12'hd08; // Dec: -760
		 575: sinewave = 12'hcfd; // Dec: -771
		 576: sinewave = 12'hcf1; // Dec: -783
		 577: sinewave = 12'hce6; // Dec: -794
		 578: sinewave = 12'hcda; // Dec: -806
		 579: sinewave = 12'hcce; // Dec: -818
		 580: sinewave = 12'hcc3; // Dec: -829
		 581: sinewave = 12'hcb8; // Dec: -840
		 582: sinewave = 12'hcac; // Dec: -852
		 583: sinewave = 12'hca1; // Dec: -863
		 584: sinewave = 12'hc95; // Dec: -875
		 585: sinewave = 12'hc8a; // Dec: -886
		 586: sinewave = 12'hc7f; // Dec: -897
		 587: sinewave = 12'hc73; // Dec: -909
		 588: sinewave = 12'hc68; // Dec: -920
		 589: sinewave = 12'hc5d; // Dec: -931
		 590: sinewave = 12'hc52; // Dec: -942
		 591: sinewave = 12'hc47; // Dec: -953
		 592: sinewave = 12'hc3c; // Dec: -964
		 593: sinewave = 12'hc30; // Dec: -976
		 594: sinewave = 12'hc25; // Dec: -987
		 595: sinewave = 12'hc1a; // Dec: -998
		 596: sinewave = 12'hc10; // Dec: -1008
		 597: sinewave = 12'hc05; // Dec: -1019
		 598: sinewave = 12'hbfa; // Dec: -1030
		 599: sinewave = 12'hbef; // Dec: -1041
		 600: sinewave = 12'hbe4; // Dec: -1052
		 601: sinewave = 12'hbd9; // Dec: -1063
		 602: sinewave = 12'hbcf; // Dec: -1073
		 603: sinewave = 12'hbc4; // Dec: -1084
		 604: sinewave = 12'hbb9; // Dec: -1095
		 605: sinewave = 12'hbaf; // Dec: -1105
		 606: sinewave = 12'hba4; // Dec: -1116
		 607: sinewave = 12'hb9a; // Dec: -1126
		 608: sinewave = 12'hb8f; // Dec: -1137
		 609: sinewave = 12'hb85; // Dec: -1147
		 610: sinewave = 12'hb7a; // Dec: -1158
		 611: sinewave = 12'hb70; // Dec: -1168
		 612: sinewave = 12'hb66; // Dec: -1178
		 613: sinewave = 12'hb5c; // Dec: -1188
		 614: sinewave = 12'hb51; // Dec: -1199
		 615: sinewave = 12'hb47; // Dec: -1209
		 616: sinewave = 12'hb3d; // Dec: -1219
		 617: sinewave = 12'hb33; // Dec: -1229
		 618: sinewave = 12'hb29; // Dec: -1239
		 619: sinewave = 12'hb1f; // Dec: -1249
		 620: sinewave = 12'hb15; // Dec: -1259
		 621: sinewave = 12'hb0b; // Dec: -1269
		 622: sinewave = 12'hb01; // Dec: -1279
		 623: sinewave = 12'haf8; // Dec: -1288
		 624: sinewave = 12'haee; // Dec: -1298
		 625: sinewave = 12'hae4; // Dec: -1308
		 626: sinewave = 12'hadb; // Dec: -1317
		 627: sinewave = 12'had1; // Dec: -1327
		 628: sinewave = 12'hac7; // Dec: -1337
		 629: sinewave = 12'habe; // Dec: -1346
		 630: sinewave = 12'hab5; // Dec: -1355
		 631: sinewave = 12'haab; // Dec: -1365
		 632: sinewave = 12'haa2; // Dec: -1374
		 633: sinewave = 12'ha99; // Dec: -1383
		 634: sinewave = 12'ha8f; // Dec: -1393
		 635: sinewave = 12'ha86; // Dec: -1402
		 636: sinewave = 12'ha7d; // Dec: -1411
		 637: sinewave = 12'ha74; // Dec: -1420
		 638: sinewave = 12'ha6b; // Dec: -1429
		 639: sinewave = 12'ha62; // Dec: -1438
		 640: sinewave = 12'ha59; // Dec: -1447
		 641: sinewave = 12'ha50; // Dec: -1456
		 642: sinewave = 12'ha47; // Dec: -1465
		 643: sinewave = 12'ha3f; // Dec: -1473
		 644: sinewave = 12'ha36; // Dec: -1482
		 645: sinewave = 12'ha2d; // Dec: -1491
		 646: sinewave = 12'ha25; // Dec: -1499
		 647: sinewave = 12'ha1c; // Dec: -1508
		 648: sinewave = 12'ha14; // Dec: -1516
		 649: sinewave = 12'ha0b; // Dec: -1525
		 650: sinewave = 12'ha03; // Dec: -1533
		 651: sinewave = 12'h9fb; // Dec: -1541
		 652: sinewave = 12'h9f2; // Dec: -1550
		 653: sinewave = 12'h9ea; // Dec: -1558
		 654: sinewave = 12'h9e2; // Dec: -1566
		 655: sinewave = 12'h9da; // Dec: -1574
		 656: sinewave = 12'h9d2; // Dec: -1582
		 657: sinewave = 12'h9ca; // Dec: -1590
		 658: sinewave = 12'h9c2; // Dec: -1598
		 659: sinewave = 12'h9bb; // Dec: -1605
		 660: sinewave = 12'h9b3; // Dec: -1613
		 661: sinewave = 12'h9ab; // Dec: -1621
		 662: sinewave = 12'h9a3; // Dec: -1629
		 663: sinewave = 12'h99c; // Dec: -1636
		 664: sinewave = 12'h994; // Dec: -1644
		 665: sinewave = 12'h98d; // Dec: -1651
		 666: sinewave = 12'h985; // Dec: -1659
		 667: sinewave = 12'h97e; // Dec: -1666
		 668: sinewave = 12'h977; // Dec: -1673
		 669: sinewave = 12'h970; // Dec: -1680
		 670: sinewave = 12'h969; // Dec: -1687
		 671: sinewave = 12'h961; // Dec: -1695
		 672: sinewave = 12'h95a; // Dec: -1702
		 673: sinewave = 12'h954; // Dec: -1708
		 674: sinewave = 12'h94d; // Dec: -1715
		 675: sinewave = 12'h946; // Dec: -1722
		 676: sinewave = 12'h93f; // Dec: -1729
		 677: sinewave = 12'h938; // Dec: -1736
		 678: sinewave = 12'h932; // Dec: -1742
		 679: sinewave = 12'h92b; // Dec: -1749
		 680: sinewave = 12'h925; // Dec: -1755
		 681: sinewave = 12'h91e; // Dec: -1762
		 682: sinewave = 12'h918; // Dec: -1768
		 683: sinewave = 12'h912; // Dec: -1774
		 684: sinewave = 12'h90b; // Dec: -1781
		 685: sinewave = 12'h905; // Dec: -1787
		 686: sinewave = 12'h8ff; // Dec: -1793
		 687: sinewave = 12'h8f9; // Dec: -1799
		 688: sinewave = 12'h8f3; // Dec: -1805
		 689: sinewave = 12'h8ed; // Dec: -1811
		 690: sinewave = 12'h8e8; // Dec: -1816
		 691: sinewave = 12'h8e2; // Dec: -1822
		 692: sinewave = 12'h8dc; // Dec: -1828
		 693: sinewave = 12'h8d6; // Dec: -1834
		 694: sinewave = 12'h8d1; // Dec: -1839
		 695: sinewave = 12'h8cb; // Dec: -1845
		 696: sinewave = 12'h8c6; // Dec: -1850
		 697: sinewave = 12'h8c1; // Dec: -1855
		 698: sinewave = 12'h8bb; // Dec: -1861
		 699: sinewave = 12'h8b6; // Dec: -1866
		 700: sinewave = 12'h8b1; // Dec: -1871
		 701: sinewave = 12'h8ac; // Dec: -1876
		 702: sinewave = 12'h8a7; // Dec: -1881
		 703: sinewave = 12'h8a2; // Dec: -1886
		 704: sinewave = 12'h89d; // Dec: -1891
		 705: sinewave = 12'h899; // Dec: -1895
		 706: sinewave = 12'h894; // Dec: -1900
		 707: sinewave = 12'h88f; // Dec: -1905
		 708: sinewave = 12'h88b; // Dec: -1909
		 709: sinewave = 12'h886; // Dec: -1914
		 710: sinewave = 12'h882; // Dec: -1918
		 711: sinewave = 12'h87d; // Dec: -1923
		 712: sinewave = 12'h879; // Dec: -1927
		 713: sinewave = 12'h875; // Dec: -1931
		 714: sinewave = 12'h871; // Dec: -1935
		 715: sinewave = 12'h86d; // Dec: -1939
		 716: sinewave = 12'h869; // Dec: -1943
		 717: sinewave = 12'h865; // Dec: -1947
		 718: sinewave = 12'h861; // Dec: -1951
		 719: sinewave = 12'h85d; // Dec: -1955
		 720: sinewave = 12'h85a; // Dec: -1958
		 721: sinewave = 12'h856; // Dec: -1962
		 722: sinewave = 12'h852; // Dec: -1966
		 723: sinewave = 12'h84f; // Dec: -1969
		 724: sinewave = 12'h84c; // Dec: -1972
		 725: sinewave = 12'h848; // Dec: -1976
		 726: sinewave = 12'h845; // Dec: -1979
		 727: sinewave = 12'h842; // Dec: -1982
		 728: sinewave = 12'h83f; // Dec: -1985
		 729: sinewave = 12'h83c; // Dec: -1988
		 730: sinewave = 12'h839; // Dec: -1991
		 731: sinewave = 12'h836; // Dec: -1994
		 732: sinewave = 12'h833; // Dec: -1997
		 733: sinewave = 12'h831; // Dec: -1999
		 734: sinewave = 12'h82e; // Dec: -2002
		 735: sinewave = 12'h82b; // Dec: -2005
		 736: sinewave = 12'h829; // Dec: -2007
		 737: sinewave = 12'h826; // Dec: -2010
		 738: sinewave = 12'h824; // Dec: -2012
		 739: sinewave = 12'h822; // Dec: -2014
		 740: sinewave = 12'h820; // Dec: -2016
		 741: sinewave = 12'h81e; // Dec: -2018
		 742: sinewave = 12'h81b; // Dec: -2021
		 743: sinewave = 12'h81a; // Dec: -2022
		 744: sinewave = 12'h818; // Dec: -2024
		 745: sinewave = 12'h816; // Dec: -2026
		 746: sinewave = 12'h814; // Dec: -2028
		 747: sinewave = 12'h812; // Dec: -2030
		 748: sinewave = 12'h811; // Dec: -2031
		 749: sinewave = 12'h80f; // Dec: -2033
		 750: sinewave = 12'h80e; // Dec: -2034
		 751: sinewave = 12'h80d; // Dec: -2035
		 752: sinewave = 12'h80b; // Dec: -2037
		 753: sinewave = 12'h80a; // Dec: -2038
		 754: sinewave = 12'h809; // Dec: -2039
		 755: sinewave = 12'h808; // Dec: -2040
		 756: sinewave = 12'h807; // Dec: -2041
		 757: sinewave = 12'h806; // Dec: -2042
		 758: sinewave = 12'h805; // Dec: -2043
		 759: sinewave = 12'h805; // Dec: -2043
		 760: sinewave = 12'h804; // Dec: -2044
		 761: sinewave = 12'h803; // Dec: -2045
		 762: sinewave = 12'h803; // Dec: -2045
		 763: sinewave = 12'h802; // Dec: -2046
		 764: sinewave = 12'h802; // Dec: -2046
		 765: sinewave = 12'h802; // Dec: -2046
		 766: sinewave = 12'h802; // Dec: -2046
		 767: sinewave = 12'h802; // Dec: -2046
		 768: sinewave = 12'h801; // Dec: -2047
		 769: sinewave = 12'h802; // Dec: -2046
		 770: sinewave = 12'h802; // Dec: -2046
		 771: sinewave = 12'h802; // Dec: -2046
		 772: sinewave = 12'h802; // Dec: -2046
		 773: sinewave = 12'h802; // Dec: -2046
		 774: sinewave = 12'h803; // Dec: -2045
		 775: sinewave = 12'h803; // Dec: -2045
		 776: sinewave = 12'h804; // Dec: -2044
		 777: sinewave = 12'h805; // Dec: -2043
		 778: sinewave = 12'h805; // Dec: -2043
		 779: sinewave = 12'h806; // Dec: -2042
		 780: sinewave = 12'h807; // Dec: -2041
		 781: sinewave = 12'h808; // Dec: -2040
		 782: sinewave = 12'h809; // Dec: -2039
		 783: sinewave = 12'h80a; // Dec: -2038
		 784: sinewave = 12'h80b; // Dec: -2037
		 785: sinewave = 12'h80d; // Dec: -2035
		 786: sinewave = 12'h80e; // Dec: -2034
		 787: sinewave = 12'h80f; // Dec: -2033
		 788: sinewave = 12'h811; // Dec: -2031
		 789: sinewave = 12'h812; // Dec: -2030
		 790: sinewave = 12'h814; // Dec: -2028
		 791: sinewave = 12'h816; // Dec: -2026
		 792: sinewave = 12'h818; // Dec: -2024
		 793: sinewave = 12'h81a; // Dec: -2022
		 794: sinewave = 12'h81b; // Dec: -2021
		 795: sinewave = 12'h81e; // Dec: -2018
		 796: sinewave = 12'h820; // Dec: -2016
		 797: sinewave = 12'h822; // Dec: -2014
		 798: sinewave = 12'h824; // Dec: -2012
		 799: sinewave = 12'h826; // Dec: -2010
		 800: sinewave = 12'h829; // Dec: -2007
		 801: sinewave = 12'h82b; // Dec: -2005
		 802: sinewave = 12'h82e; // Dec: -2002
		 803: sinewave = 12'h831; // Dec: -1999
		 804: sinewave = 12'h833; // Dec: -1997
		 805: sinewave = 12'h836; // Dec: -1994
		 806: sinewave = 12'h839; // Dec: -1991
		 807: sinewave = 12'h83c; // Dec: -1988
		 808: sinewave = 12'h83f; // Dec: -1985
		 809: sinewave = 12'h842; // Dec: -1982
		 810: sinewave = 12'h845; // Dec: -1979
		 811: sinewave = 12'h848; // Dec: -1976
		 812: sinewave = 12'h84c; // Dec: -1972
		 813: sinewave = 12'h84f; // Dec: -1969
		 814: sinewave = 12'h852; // Dec: -1966
		 815: sinewave = 12'h856; // Dec: -1962
		 816: sinewave = 12'h85a; // Dec: -1958
		 817: sinewave = 12'h85d; // Dec: -1955
		 818: sinewave = 12'h861; // Dec: -1951
		 819: sinewave = 12'h865; // Dec: -1947
		 820: sinewave = 12'h869; // Dec: -1943
		 821: sinewave = 12'h86d; // Dec: -1939
		 822: sinewave = 12'h871; // Dec: -1935
		 823: sinewave = 12'h875; // Dec: -1931
		 824: sinewave = 12'h879; // Dec: -1927
		 825: sinewave = 12'h87d; // Dec: -1923
		 826: sinewave = 12'h882; // Dec: -1918
		 827: sinewave = 12'h886; // Dec: -1914
		 828: sinewave = 12'h88b; // Dec: -1909
		 829: sinewave = 12'h88f; // Dec: -1905
		 830: sinewave = 12'h894; // Dec: -1900
		 831: sinewave = 12'h899; // Dec: -1895
		 832: sinewave = 12'h89d; // Dec: -1891
		 833: sinewave = 12'h8a2; // Dec: -1886
		 834: sinewave = 12'h8a7; // Dec: -1881
		 835: sinewave = 12'h8ac; // Dec: -1876
		 836: sinewave = 12'h8b1; // Dec: -1871
		 837: sinewave = 12'h8b6; // Dec: -1866
		 838: sinewave = 12'h8bb; // Dec: -1861
		 839: sinewave = 12'h8c1; // Dec: -1855
		 840: sinewave = 12'h8c6; // Dec: -1850
		 841: sinewave = 12'h8cb; // Dec: -1845
		 842: sinewave = 12'h8d1; // Dec: -1839
		 843: sinewave = 12'h8d6; // Dec: -1834
		 844: sinewave = 12'h8dc; // Dec: -1828
		 845: sinewave = 12'h8e2; // Dec: -1822
		 846: sinewave = 12'h8e8; // Dec: -1816
		 847: sinewave = 12'h8ed; // Dec: -1811
		 848: sinewave = 12'h8f3; // Dec: -1805
		 849: sinewave = 12'h8f9; // Dec: -1799
		 850: sinewave = 12'h8ff; // Dec: -1793
		 851: sinewave = 12'h905; // Dec: -1787
		 852: sinewave = 12'h90b; // Dec: -1781
		 853: sinewave = 12'h912; // Dec: -1774
		 854: sinewave = 12'h918; // Dec: -1768
		 855: sinewave = 12'h91e; // Dec: -1762
		 856: sinewave = 12'h925; // Dec: -1755
		 857: sinewave = 12'h92b; // Dec: -1749
		 858: sinewave = 12'h932; // Dec: -1742
		 859: sinewave = 12'h938; // Dec: -1736
		 860: sinewave = 12'h93f; // Dec: -1729
		 861: sinewave = 12'h946; // Dec: -1722
		 862: sinewave = 12'h94d; // Dec: -1715
		 863: sinewave = 12'h954; // Dec: -1708
		 864: sinewave = 12'h95a; // Dec: -1702
		 865: sinewave = 12'h961; // Dec: -1695
		 866: sinewave = 12'h969; // Dec: -1687
		 867: sinewave = 12'h970; // Dec: -1680
		 868: sinewave = 12'h977; // Dec: -1673
		 869: sinewave = 12'h97e; // Dec: -1666
		 870: sinewave = 12'h985; // Dec: -1659
		 871: sinewave = 12'h98d; // Dec: -1651
		 872: sinewave = 12'h994; // Dec: -1644
		 873: sinewave = 12'h99c; // Dec: -1636
		 874: sinewave = 12'h9a3; // Dec: -1629
		 875: sinewave = 12'h9ab; // Dec: -1621
		 876: sinewave = 12'h9b3; // Dec: -1613
		 877: sinewave = 12'h9bb; // Dec: -1605
		 878: sinewave = 12'h9c2; // Dec: -1598
		 879: sinewave = 12'h9ca; // Dec: -1590
		 880: sinewave = 12'h9d2; // Dec: -1582
		 881: sinewave = 12'h9da; // Dec: -1574
		 882: sinewave = 12'h9e2; // Dec: -1566
		 883: sinewave = 12'h9ea; // Dec: -1558
		 884: sinewave = 12'h9f2; // Dec: -1550
		 885: sinewave = 12'h9fb; // Dec: -1541
		 886: sinewave = 12'ha03; // Dec: -1533
		 887: sinewave = 12'ha0b; // Dec: -1525
		 888: sinewave = 12'ha14; // Dec: -1516
		 889: sinewave = 12'ha1c; // Dec: -1508
		 890: sinewave = 12'ha25; // Dec: -1499
		 891: sinewave = 12'ha2d; // Dec: -1491
		 892: sinewave = 12'ha36; // Dec: -1482
		 893: sinewave = 12'ha3f; // Dec: -1473
		 894: sinewave = 12'ha47; // Dec: -1465
		 895: sinewave = 12'ha50; // Dec: -1456
		 896: sinewave = 12'ha59; // Dec: -1447
		 897: sinewave = 12'ha62; // Dec: -1438
		 898: sinewave = 12'ha6b; // Dec: -1429
		 899: sinewave = 12'ha74; // Dec: -1420
		 900: sinewave = 12'ha7d; // Dec: -1411
		 901: sinewave = 12'ha86; // Dec: -1402
		 902: sinewave = 12'ha8f; // Dec: -1393
		 903: sinewave = 12'ha99; // Dec: -1383
		 904: sinewave = 12'haa2; // Dec: -1374
		 905: sinewave = 12'haab; // Dec: -1365
		 906: sinewave = 12'hab5; // Dec: -1355
		 907: sinewave = 12'habe; // Dec: -1346
		 908: sinewave = 12'hac7; // Dec: -1337
		 909: sinewave = 12'had1; // Dec: -1327
		 910: sinewave = 12'hadb; // Dec: -1317
		 911: sinewave = 12'hae4; // Dec: -1308
		 912: sinewave = 12'haee; // Dec: -1298
		 913: sinewave = 12'haf8; // Dec: -1288
		 914: sinewave = 12'hb01; // Dec: -1279
		 915: sinewave = 12'hb0b; // Dec: -1269
		 916: sinewave = 12'hb15; // Dec: -1259
		 917: sinewave = 12'hb1f; // Dec: -1249
		 918: sinewave = 12'hb29; // Dec: -1239
		 919: sinewave = 12'hb33; // Dec: -1229
		 920: sinewave = 12'hb3d; // Dec: -1219
		 921: sinewave = 12'hb47; // Dec: -1209
		 922: sinewave = 12'hb51; // Dec: -1199
		 923: sinewave = 12'hb5c; // Dec: -1188
		 924: sinewave = 12'hb66; // Dec: -1178
		 925: sinewave = 12'hb70; // Dec: -1168
		 926: sinewave = 12'hb7a; // Dec: -1158
		 927: sinewave = 12'hb85; // Dec: -1147
		 928: sinewave = 12'hb8f; // Dec: -1137
		 929: sinewave = 12'hb9a; // Dec: -1126
		 930: sinewave = 12'hba4; // Dec: -1116
		 931: sinewave = 12'hbaf; // Dec: -1105
		 932: sinewave = 12'hbb9; // Dec: -1095
		 933: sinewave = 12'hbc4; // Dec: -1084
		 934: sinewave = 12'hbcf; // Dec: -1073
		 935: sinewave = 12'hbd9; // Dec: -1063
		 936: sinewave = 12'hbe4; // Dec: -1052
		 937: sinewave = 12'hbef; // Dec: -1041
		 938: sinewave = 12'hbfa; // Dec: -1030
		 939: sinewave = 12'hc05; // Dec: -1019
		 940: sinewave = 12'hc10; // Dec: -1008
		 941: sinewave = 12'hc1a; // Dec: -998
		 942: sinewave = 12'hc25; // Dec: -987
		 943: sinewave = 12'hc30; // Dec: -976
		 944: sinewave = 12'hc3c; // Dec: -964
		 945: sinewave = 12'hc47; // Dec: -953
		 946: sinewave = 12'hc52; // Dec: -942
		 947: sinewave = 12'hc5d; // Dec: -931
		 948: sinewave = 12'hc68; // Dec: -920
		 949: sinewave = 12'hc73; // Dec: -909
		 950: sinewave = 12'hc7f; // Dec: -897
		 951: sinewave = 12'hc8a; // Dec: -886
		 952: sinewave = 12'hc95; // Dec: -875
		 953: sinewave = 12'hca1; // Dec: -863
		 954: sinewave = 12'hcac; // Dec: -852
		 955: sinewave = 12'hcb8; // Dec: -840
		 956: sinewave = 12'hcc3; // Dec: -829
		 957: sinewave = 12'hcce; // Dec: -818
		 958: sinewave = 12'hcda; // Dec: -806
		 959: sinewave = 12'hce6; // Dec: -794
		 960: sinewave = 12'hcf1; // Dec: -783
		 961: sinewave = 12'hcfd; // Dec: -771
		 962: sinewave = 12'hd08; // Dec: -760
		 963: sinewave = 12'hd14; // Dec: -748
		 964: sinewave = 12'hd20; // Dec: -736
		 965: sinewave = 12'hd2c; // Dec: -724
		 966: sinewave = 12'hd37; // Dec: -713
		 967: sinewave = 12'hd43; // Dec: -701
		 968: sinewave = 12'hd4f; // Dec: -689
		 969: sinewave = 12'hd5b; // Dec: -677
		 970: sinewave = 12'hd67; // Dec: -665
		 971: sinewave = 12'hd72; // Dec: -654
		 972: sinewave = 12'hd7e; // Dec: -642
		 973: sinewave = 12'hd8a; // Dec: -630
		 974: sinewave = 12'hd96; // Dec: -618
		 975: sinewave = 12'hda2; // Dec: -606
		 976: sinewave = 12'hdae; // Dec: -594
		 977: sinewave = 12'hdba; // Dec: -582
		 978: sinewave = 12'hdc6; // Dec: -570
		 979: sinewave = 12'hdd2; // Dec: -558
		 980: sinewave = 12'hddf; // Dec: -545
		 981: sinewave = 12'hdeb; // Dec: -533
		 982: sinewave = 12'hdf7; // Dec: -521
		 983: sinewave = 12'he03; // Dec: -509
		 984: sinewave = 12'he0f; // Dec: -497
		 985: sinewave = 12'he1b; // Dec: -485
		 986: sinewave = 12'he28; // Dec: -472
		 987: sinewave = 12'he34; // Dec: -460
		 988: sinewave = 12'he40; // Dec: -448
		 989: sinewave = 12'he4c; // Dec: -436
		 990: sinewave = 12'he59; // Dec: -423
		 991: sinewave = 12'he65; // Dec: -411
		 992: sinewave = 12'he71; // Dec: -399
		 993: sinewave = 12'he7d; // Dec: -387
		 994: sinewave = 12'he8a; // Dec: -374
		 995: sinewave = 12'he96; // Dec: -362
		 996: sinewave = 12'hea3; // Dec: -349
		 997: sinewave = 12'heaf; // Dec: -337
		 998: sinewave = 12'hebb; // Dec: -325
		 999: sinewave = 12'hec8; // Dec: -312
		1000: sinewave = 12'hed4; // Dec: -300
		1001: sinewave = 12'hee1; // Dec: -287
		1002: sinewave = 12'heed; // Dec: -275
		1003: sinewave = 12'hef9; // Dec: -263
		1004: sinewave = 12'hf06; // Dec: -250
		1005: sinewave = 12'hf12; // Dec: -238
		1006: sinewave = 12'hf1f; // Dec: -225
		1007: sinewave = 12'hf2b; // Dec: -213
		1008: sinewave = 12'hf38; // Dec: -200
		1009: sinewave = 12'hf44; // Dec: -188
		1010: sinewave = 12'hf51; // Dec: -175
		1011: sinewave = 12'hf5d; // Dec: -163
		1012: sinewave = 12'hf6a; // Dec: -150
		1013: sinewave = 12'hf76; // Dec: -138
		1014: sinewave = 12'hf83; // Dec: -125
		1015: sinewave = 12'hf90; // Dec: -112
		1016: sinewave = 12'hf9c; // Dec: -100
		1017: sinewave = 12'hfa9; // Dec: -87
		1018: sinewave = 12'hfb5; // Dec: -75
		1019: sinewave = 12'hfc2; // Dec: -62
		1020: sinewave = 12'hfce; // Dec: -50
		1021: sinewave = 12'hfdb; // Dec: -37
		1022: sinewave = 12'hfe7; // Dec: -25
		1023: sinewave = 12'hff4; // Dec: -12
		endcase

end

endmodule
