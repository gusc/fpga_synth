`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Tomass Lacis
// 
// Create Date:    16:14:10 05/19/2018 
// Design Name: 
// Module Name:    SampleGenerator 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SampleGenerator(
	inCLK,
	inWaveMode,
	inSampleClockCE,
	inMidiFrequencyIndex,	
	outSample
);
	// SOURCES USED: 
	// 1. http://zipcpu.com/dsp/2017/07/11/simplest-sinewave-generator.html
	
	// === PARAMETERS ===
	parameter SAMPLE_CLOCK_RATE_HZ = 44100;
	parameter N = 32; // Phase bit width
	parameter M = 12; // Sample output bit width
	
	// === I/O ===
	input inCLK;
	input [1:0] inWaveMode;
	input inSampleClockCE;
	input [6:0] inMidiFrequencyIndex;
	output reg [M-1:0] outSample;
	
	// === REGISTERS ===
	reg [N-1:0] phase = 0; // 32bit phase
	
	// === FREQUENCY STEP TABLE ==
	reg [N-1:0] frequency_step [127:0];
	initial begin
		// Formula for frequency step: (2^N * FREQ_Z) / SAMPLE_CLOCK_RATE_HZ
		frequency_step[0]   = 796175910;
		frequency_step[1]   = 843508202;
		frequency_step[2]   = 893762242;
		frequency_step[3]   = 946840636;
		frequency_step[4]   = 1003132951;
		frequency_step[5]   = 1062833970;
		frequency_step[6]   = 1126041085;
		frequency_step[7]   = 1192949079;
		frequency_step[8]   = 1263947518;
		frequency_step[9]   = 1339133794;
		frequency_step[10]  = 1418702689;
		frequency_step[11]  = 1503043770;
		frequency_step[12]  = 1592449212;
		frequency_step[13]  = 1687113797;
		frequency_step[14]  = 1787524484;
		frequency_step[15]  = 1893778663;
		frequency_step[16]  = 2006363293;
		frequency_step[17]  = 2125667941;
		frequency_step[18]  = 2252082171;
		frequency_step[19]  = 2385995550;
		frequency_step[20]  = 2527895037;
		frequency_step[21]  = 2678267588;
		frequency_step[22]  = 2837502770;
		frequency_step[23]  = 3006184932;
		frequency_step[24]  = 3184995815;
		frequency_step[25]  = 3374324986;
		frequency_step[26]  = 3575048968;
		frequency_step[27]  = 3787557327;
		frequency_step[28]  = 4012823979;
		frequency_step[29]  = 4251433273;
		frequency_step[30]  = 209294438;
		frequency_step[31]  = 477121196;
		frequency_step[32]  = 760920169;
		frequency_step[33]  = 1061567880;
		frequency_step[34]  = 1380038244;
		frequency_step[35]  = 1717499960;
		frequency_step[36]  = 2075024335;
		frequency_step[37]  = 2453780068;
		frequency_step[38]  = 2855130640;
		frequency_step[39]  = 3280244750;
		frequency_step[40]  = 3730680663;
		frequency_step[41]  = 4207996643;
		frequency_step[42]  = 418588876;
		frequency_step[43]  = 954242393;
		frequency_step[44]  = 1521840339;
		frequency_step[45]  = 2123135760;
		frequency_step[46]  = 2760076489;
		frequency_step[47]  = 3434999921;
		frequency_step[48]  = 4150048671;
		frequency_step[49]  = 612690232;
		frequency_step[50]  = 1415293985;
		frequency_step[51]  = 2265619596;
		frequency_step[52]  = 3166491421;
		frequency_step[53]  = 4121025990;
		frequency_step[54]  = 837275143;
		frequency_step[55]  = 1908582179;
		frequency_step[56]  = 3043680678;
		frequency_step[57]  = 4246271521;
		frequency_step[58]  = 1225283073;
		frequency_step[59]  = 2575129938;
		frequency_step[60]  = 4005227438;
		frequency_step[61]  = 1225380465;
		frequency_step[62]  = 2830587970;
		frequency_step[63]  = 236271897;
		frequency_step[64]  = 2038112938;
		frequency_step[65]  = 3947084684;
		frequency_step[66]  = 1674550287;
		frequency_step[67]  = 3817261749;
		frequency_step[68]  = 1792394061;
		frequency_step[69]  = 4197575747;
		frequency_step[70]  = 2450663538;
		frequency_step[71]  = 855389971;
		frequency_step[72]  = 3715584973;
		frequency_step[73]  = 2450858322;
		frequency_step[74]  = 1366306036;
		frequency_step[75]  = 472641185;
		frequency_step[76]  = 4076323269;
		frequency_step[77]  = 3599202072;
		frequency_step[78]  = 3349100575;
		frequency_step[79]  = 3339556203;
		frequency_step[80]  = 3584885514;
		frequency_step[81]  = 4100184198;
		frequency_step[82]  = 606457173;
		frequency_step[83]  = 1710779943;
		frequency_step[84]  = 3136202650;
		frequency_step[85]  = 606749348;
		frequency_step[86]  = 2732709463;
		frequency_step[87]  = 945379762;
		frequency_step[88]  = 3857679242;
		frequency_step[89]  = 2903436848;
		frequency_step[90]  = 2403331246;
		frequency_step[91]  = 2384242502;
		frequency_step[92]  = 2874803733;
		frequency_step[93]  = 3905401101;
		frequency_step[94]  = 1213011738;
		frequency_step[95]  = 3421657279;
		frequency_step[96]  = 1977438004;
		frequency_step[97]  = 1213596087;
		frequency_step[98]  = 1170451631;
		frequency_step[99]  = 1890856917;
		frequency_step[100] = 3420391189;
		frequency_step[101] = 1512003792;
		frequency_step[102] = 511792588;
		frequency_step[103] = 473615101;
		frequency_step[104] = 1454737562;
		frequency_step[105] = 3515834906;
		frequency_step[106] = 2426023477;
		frequency_step[107] = 2548347262;
		frequency_step[108] = 3954973399;
		frequency_step[109] = 2427192175;
		frequency_step[110] = 2340903263;
		frequency_step[111] = 3781811226;
		frequency_step[112] = 2545815082;
		frequency_step[113] = 3024104977;
		frequency_step[114] = 1023585176;
		frequency_step[115] = 947230202;
		frequency_step[116] = 2909572516;
		frequency_step[117] = 2736702517;
		frequency_step[118] = 557079658;
		frequency_step[119] = 801727228;
		frequency_step[120] = 3614979503;
		frequency_step[121] = 559417055;
		frequency_step[122] = 386839231;
		frequency_step[123] = 3268752547;
		frequency_step[124] = 796760259;
		frequency_step[125] = 1753340050;
		frequency_step[126] = 2047267744;
		frequency_step[127] = 1894557796;
	end
	
	// === SINEWAVE TABLE (from 8-top-bit phase) ==
	reg [M-1:0] sinewave [1023:0];
	initial begin
		sinewave[0] = 12'h00;
		sinewave[1] = 12'h0c;
		sinewave[2] = 12'h19;
		sinewave[3] = 12'h25;
		sinewave[4] = 12'h32;
		sinewave[5] = 12'h3e;
		sinewave[6] = 12'h4b;
		sinewave[7] = 12'h57;
		sinewave[8] = 12'h64;
		sinewave[9] = 12'h70;
		sinewave[10] = 12'h7d;
		sinewave[11] = 12'h8a;
		sinewave[12] = 12'h96;
		sinewave[13] = 12'ha3;
		sinewave[14] = 12'haf;
		sinewave[15] = 12'hbc;
		sinewave[16] = 12'hc8;
		sinewave[17] = 12'hd5;
		sinewave[18] = 12'he1;
		sinewave[19] = 12'hee;
		sinewave[20] = 12'hfa;
		sinewave[21] = 12'h107;
		sinewave[22] = 12'h113;
		sinewave[23] = 12'h11f;
		sinewave[24] = 12'h12c;
		sinewave[25] = 12'h138;
		sinewave[26] = 12'h145;
		sinewave[27] = 12'h151;
		sinewave[28] = 12'h15d;
		sinewave[29] = 12'h16a;
		sinewave[30] = 12'h176;
		sinewave[31] = 12'h183;
		sinewave[32] = 12'h18f;
		sinewave[33] = 12'h19b;
		sinewave[34] = 12'h1a7;
		sinewave[35] = 12'h1b4;
		sinewave[36] = 12'h1c0;
		sinewave[37] = 12'h1cc;
		sinewave[38] = 12'h1d8;
		sinewave[39] = 12'h1e5;
		sinewave[40] = 12'h1f1;
		sinewave[41] = 12'h1fd;
		sinewave[42] = 12'h209;
		sinewave[43] = 12'h215;
		sinewave[44] = 12'h221;
		sinewave[45] = 12'h22e;
		sinewave[46] = 12'h23a;
		sinewave[47] = 12'h246;
		sinewave[48] = 12'h252;
		sinewave[49] = 12'h25e;
		sinewave[50] = 12'h26a;
		sinewave[51] = 12'h276;
		sinewave[52] = 12'h282;
		sinewave[53] = 12'h28e;
		sinewave[54] = 12'h299;
		sinewave[55] = 12'h2a5;
		sinewave[56] = 12'h2b1;
		sinewave[57] = 12'h2bd;
		sinewave[58] = 12'h2c9;
		sinewave[59] = 12'h2d4;
		sinewave[60] = 12'h2e0;
		sinewave[61] = 12'h2ec;
		sinewave[62] = 12'h2f8;
		sinewave[63] = 12'h303;
		sinewave[64] = 12'h30f;
		sinewave[65] = 12'h31a;
		sinewave[66] = 12'h326;
		sinewave[67] = 12'h332;
		sinewave[68] = 12'h33d;
		sinewave[69] = 12'h348;
		sinewave[70] = 12'h354;
		sinewave[71] = 12'h35f;
		sinewave[72] = 12'h36b;
		sinewave[73] = 12'h376;
		sinewave[74] = 12'h381;
		sinewave[75] = 12'h38d;
		sinewave[76] = 12'h398;
		sinewave[77] = 12'h3a3;
		sinewave[78] = 12'h3ae;
		sinewave[79] = 12'h3b9;
		sinewave[80] = 12'h3c4;
		sinewave[81] = 12'h3d0;
		sinewave[82] = 12'h3db;
		sinewave[83] = 12'h3e6;
		sinewave[84] = 12'h3f0;
		sinewave[85] = 12'h3fb;
		sinewave[86] = 12'h406;
		sinewave[87] = 12'h411;
		sinewave[88] = 12'h41c;
		sinewave[89] = 12'h427;
		sinewave[90] = 12'h431;
		sinewave[91] = 12'h43c;
		sinewave[92] = 12'h447;
		sinewave[93] = 12'h451;
		sinewave[94] = 12'h45c;
		sinewave[95] = 12'h466;
		sinewave[96] = 12'h471;
		sinewave[97] = 12'h47b;
		sinewave[98] = 12'h486;
		sinewave[99] = 12'h490;
		sinewave[100] = 12'h49a;
		sinewave[101] = 12'h4a4;
		sinewave[102] = 12'h4af;
		sinewave[103] = 12'h4b9;
		sinewave[104] = 12'h4c3;
		sinewave[105] = 12'h4cd;
		sinewave[106] = 12'h4d7;
		sinewave[107] = 12'h4e1;
		sinewave[108] = 12'h4eb;
		sinewave[109] = 12'h4f5;
		sinewave[110] = 12'h4ff;
		sinewave[111] = 12'h508;
		sinewave[112] = 12'h512;
		sinewave[113] = 12'h51c;
		sinewave[114] = 12'h525;
		sinewave[115] = 12'h52f;
		sinewave[116] = 12'h539;
		sinewave[117] = 12'h542;
		sinewave[118] = 12'h54b;
		sinewave[119] = 12'h555;
		sinewave[120] = 12'h55e;
		sinewave[121] = 12'h567;
		sinewave[122] = 12'h571;
		sinewave[123] = 12'h57a;
		sinewave[124] = 12'h583;
		sinewave[125] = 12'h58c;
		sinewave[126] = 12'h595;
		sinewave[127] = 12'h59e;
		sinewave[128] = 12'h5a7;
		sinewave[129] = 12'h5b0;
		sinewave[130] = 12'h5b9;
		sinewave[131] = 12'h5c1;
		sinewave[132] = 12'h5ca;
		sinewave[133] = 12'h5d3;
		sinewave[134] = 12'h5db;
		sinewave[135] = 12'h5e4;
		sinewave[136] = 12'h5ec;
		sinewave[137] = 12'h5f5;
		sinewave[138] = 12'h5fd;
		sinewave[139] = 12'h605;
		sinewave[140] = 12'h60e;
		sinewave[141] = 12'h616;
		sinewave[142] = 12'h61e;
		sinewave[143] = 12'h626;
		sinewave[144] = 12'h62e;
		sinewave[145] = 12'h636;
		sinewave[146] = 12'h63e;
		sinewave[147] = 12'h645;
		sinewave[148] = 12'h64d;
		sinewave[149] = 12'h655;
		sinewave[150] = 12'h65d;
		sinewave[151] = 12'h664;
		sinewave[152] = 12'h66c;
		sinewave[153] = 12'h673;
		sinewave[154] = 12'h67b;
		sinewave[155] = 12'h682;
		sinewave[156] = 12'h689;
		sinewave[157] = 12'h690;
		sinewave[158] = 12'h697;
		sinewave[159] = 12'h69f;
		sinewave[160] = 12'h6a6;
		sinewave[161] = 12'h6ac;
		sinewave[162] = 12'h6b3;
		sinewave[163] = 12'h6ba;
		sinewave[164] = 12'h6c1;
		sinewave[165] = 12'h6c8;
		sinewave[166] = 12'h6ce;
		sinewave[167] = 12'h6d5;
		sinewave[168] = 12'h6db;
		sinewave[169] = 12'h6e2;
		sinewave[170] = 12'h6e8;
		sinewave[171] = 12'h6ee;
		sinewave[172] = 12'h6f5;
		sinewave[173] = 12'h6fb;
		sinewave[174] = 12'h701;
		sinewave[175] = 12'h707;
		sinewave[176] = 12'h70d;
		sinewave[177] = 12'h713;
		sinewave[178] = 12'h718;
		sinewave[179] = 12'h71e;
		sinewave[180] = 12'h724;
		sinewave[181] = 12'h72a;
		sinewave[182] = 12'h72f;
		sinewave[183] = 12'h735;
		sinewave[184] = 12'h73a;
		sinewave[185] = 12'h73f;
		sinewave[186] = 12'h745;
		sinewave[187] = 12'h74a;
		sinewave[188] = 12'h74f;
		sinewave[189] = 12'h754;
		sinewave[190] = 12'h759;
		sinewave[191] = 12'h75e;
		sinewave[192] = 12'h763;
		sinewave[193] = 12'h767;
		sinewave[194] = 12'h76c;
		sinewave[195] = 12'h771;
		sinewave[196] = 12'h775;
		sinewave[197] = 12'h77a;
		sinewave[198] = 12'h77e;
		sinewave[199] = 12'h783;
		sinewave[200] = 12'h787;
		sinewave[201] = 12'h78b;
		sinewave[202] = 12'h78f;
		sinewave[203] = 12'h793;
		sinewave[204] = 12'h797;
		sinewave[205] = 12'h79b;
		sinewave[206] = 12'h79f;
		sinewave[207] = 12'h7a3;
		sinewave[208] = 12'h7a6;
		sinewave[209] = 12'h7aa;
		sinewave[210] = 12'h7ae;
		sinewave[211] = 12'h7b1;
		sinewave[212] = 12'h7b4;
		sinewave[213] = 12'h7b8;
		sinewave[214] = 12'h7bb;
		sinewave[215] = 12'h7be;
		sinewave[216] = 12'h7c1;
		sinewave[217] = 12'h7c4;
		sinewave[218] = 12'h7c7;
		sinewave[219] = 12'h7ca;
		sinewave[220] = 12'h7cd;
		sinewave[221] = 12'h7cf;
		sinewave[222] = 12'h7d2;
		sinewave[223] = 12'h7d5;
		sinewave[224] = 12'h7d7;
		sinewave[225] = 12'h7da;
		sinewave[226] = 12'h7dc;
		sinewave[227] = 12'h7de;
		sinewave[228] = 12'h7e0;
		sinewave[229] = 12'h7e2;
		sinewave[230] = 12'h7e5;
		sinewave[231] = 12'h7e6;
		sinewave[232] = 12'h7e8;
		sinewave[233] = 12'h7ea;
		sinewave[234] = 12'h7ec;
		sinewave[235] = 12'h7ee;
		sinewave[236] = 12'h7ef;
		sinewave[237] = 12'h7f1;
		sinewave[238] = 12'h7f2;
		sinewave[239] = 12'h7f3;
		sinewave[240] = 12'h7f5;
		sinewave[241] = 12'h7f6;
		sinewave[242] = 12'h7f7;
		sinewave[243] = 12'h7f8;
		sinewave[244] = 12'h7f9;
		sinewave[245] = 12'h7fa;
		sinewave[246] = 12'h7fb;
		sinewave[247] = 12'h7fb;
		sinewave[248] = 12'h7fc;
		sinewave[249] = 12'h7fd;
		sinewave[250] = 12'h7fd;
		sinewave[251] = 12'h7fe;
		sinewave[252] = 12'h7fe;
		sinewave[253] = 12'h7fe;
		sinewave[254] = 12'h7fe;
		sinewave[255] = 12'h7fe;
		sinewave[256] = 12'h7ff;
		sinewave[257] = 12'h7fe;
		sinewave[258] = 12'h7fe;
		sinewave[259] = 12'h7fe;
		sinewave[260] = 12'h7fe;
		sinewave[261] = 12'h7fe;
		sinewave[262] = 12'h7fd;
		sinewave[263] = 12'h7fd;
		sinewave[264] = 12'h7fc;
		sinewave[265] = 12'h7fb;
		sinewave[266] = 12'h7fb;
		sinewave[267] = 12'h7fa;
		sinewave[268] = 12'h7f9;
		sinewave[269] = 12'h7f8;
		sinewave[270] = 12'h7f7;
		sinewave[271] = 12'h7f6;
		sinewave[272] = 12'h7f5;
		sinewave[273] = 12'h7f3;
		sinewave[274] = 12'h7f2;
		sinewave[275] = 12'h7f1;
		sinewave[276] = 12'h7ef;
		sinewave[277] = 12'h7ee;
		sinewave[278] = 12'h7ec;
		sinewave[279] = 12'h7ea;
		sinewave[280] = 12'h7e8;
		sinewave[281] = 12'h7e6;
		sinewave[282] = 12'h7e5;
		sinewave[283] = 12'h7e2;
		sinewave[284] = 12'h7e0;
		sinewave[285] = 12'h7de;
		sinewave[286] = 12'h7dc;
		sinewave[287] = 12'h7da;
		sinewave[288] = 12'h7d7;
		sinewave[289] = 12'h7d5;
		sinewave[290] = 12'h7d2;
		sinewave[291] = 12'h7cf;
		sinewave[292] = 12'h7cd;
		sinewave[293] = 12'h7ca;
		sinewave[294] = 12'h7c7;
		sinewave[295] = 12'h7c4;
		sinewave[296] = 12'h7c1;
		sinewave[297] = 12'h7be;
		sinewave[298] = 12'h7bb;
		sinewave[299] = 12'h7b8;
		sinewave[300] = 12'h7b4;
		sinewave[301] = 12'h7b1;
		sinewave[302] = 12'h7ae;
		sinewave[303] = 12'h7aa;
		sinewave[304] = 12'h7a6;
		sinewave[305] = 12'h7a3;
		sinewave[306] = 12'h79f;
		sinewave[307] = 12'h79b;
		sinewave[308] = 12'h797;
		sinewave[309] = 12'h793;
		sinewave[310] = 12'h78f;
		sinewave[311] = 12'h78b;
		sinewave[312] = 12'h787;
		sinewave[313] = 12'h783;
		sinewave[314] = 12'h77e;
		sinewave[315] = 12'h77a;
		sinewave[316] = 12'h775;
		sinewave[317] = 12'h771;
		sinewave[318] = 12'h76c;
		sinewave[319] = 12'h767;
		sinewave[320] = 12'h763;
		sinewave[321] = 12'h75e;
		sinewave[322] = 12'h759;
		sinewave[323] = 12'h754;
		sinewave[324] = 12'h74f;
		sinewave[325] = 12'h74a;
		sinewave[326] = 12'h745;
		sinewave[327] = 12'h73f;
		sinewave[328] = 12'h73a;
		sinewave[329] = 12'h735;
		sinewave[330] = 12'h72f;
		sinewave[331] = 12'h72a;
		sinewave[332] = 12'h724;
		sinewave[333] = 12'h71e;
		sinewave[334] = 12'h718;
		sinewave[335] = 12'h713;
		sinewave[336] = 12'h70d;
		sinewave[337] = 12'h707;
		sinewave[338] = 12'h701;
		sinewave[339] = 12'h6fb;
		sinewave[340] = 12'h6f5;
		sinewave[341] = 12'h6ee;
		sinewave[342] = 12'h6e8;
		sinewave[343] = 12'h6e2;
		sinewave[344] = 12'h6db;
		sinewave[345] = 12'h6d5;
		sinewave[346] = 12'h6ce;
		sinewave[347] = 12'h6c8;
		sinewave[348] = 12'h6c1;
		sinewave[349] = 12'h6ba;
		sinewave[350] = 12'h6b3;
		sinewave[351] = 12'h6ac;
		sinewave[352] = 12'h6a6;
		sinewave[353] = 12'h69f;
		sinewave[354] = 12'h697;
		sinewave[355] = 12'h690;
		sinewave[356] = 12'h689;
		sinewave[357] = 12'h682;
		sinewave[358] = 12'h67b;
		sinewave[359] = 12'h673;
		sinewave[360] = 12'h66c;
		sinewave[361] = 12'h664;
		sinewave[362] = 12'h65d;
		sinewave[363] = 12'h655;
		sinewave[364] = 12'h64d;
		sinewave[365] = 12'h645;
		sinewave[366] = 12'h63e;
		sinewave[367] = 12'h636;
		sinewave[368] = 12'h62e;
		sinewave[369] = 12'h626;
		sinewave[370] = 12'h61e;
		sinewave[371] = 12'h616;
		sinewave[372] = 12'h60e;
		sinewave[373] = 12'h605;
		sinewave[374] = 12'h5fd;
		sinewave[375] = 12'h5f5;
		sinewave[376] = 12'h5ec;
		sinewave[377] = 12'h5e4;
		sinewave[378] = 12'h5db;
		sinewave[379] = 12'h5d3;
		sinewave[380] = 12'h5ca;
		sinewave[381] = 12'h5c1;
		sinewave[382] = 12'h5b9;
		sinewave[383] = 12'h5b0;
		sinewave[384] = 12'h5a7;
		sinewave[385] = 12'h59e;
		sinewave[386] = 12'h595;
		sinewave[387] = 12'h58c;
		sinewave[388] = 12'h583;
		sinewave[389] = 12'h57a;
		sinewave[390] = 12'h571;
		sinewave[391] = 12'h567;
		sinewave[392] = 12'h55e;
		sinewave[393] = 12'h555;
		sinewave[394] = 12'h54b;
		sinewave[395] = 12'h542;
		sinewave[396] = 12'h539;
		sinewave[397] = 12'h52f;
		sinewave[398] = 12'h525;
		sinewave[399] = 12'h51c;
		sinewave[400] = 12'h512;
		sinewave[401] = 12'h508;
		sinewave[402] = 12'h4ff;
		sinewave[403] = 12'h4f5;
		sinewave[404] = 12'h4eb;
		sinewave[405] = 12'h4e1;
		sinewave[406] = 12'h4d7;
		sinewave[407] = 12'h4cd;
		sinewave[408] = 12'h4c3;
		sinewave[409] = 12'h4b9;
		sinewave[410] = 12'h4af;
		sinewave[411] = 12'h4a4;
		sinewave[412] = 12'h49a;
		sinewave[413] = 12'h490;
		sinewave[414] = 12'h486;
		sinewave[415] = 12'h47b;
		sinewave[416] = 12'h471;
		sinewave[417] = 12'h466;
		sinewave[418] = 12'h45c;
		sinewave[419] = 12'h451;
		sinewave[420] = 12'h447;
		sinewave[421] = 12'h43c;
		sinewave[422] = 12'h431;
		sinewave[423] = 12'h427;
		sinewave[424] = 12'h41c;
		sinewave[425] = 12'h411;
		sinewave[426] = 12'h406;
		sinewave[427] = 12'h3fb;
		sinewave[428] = 12'h3f0;
		sinewave[429] = 12'h3e6;
		sinewave[430] = 12'h3db;
		sinewave[431] = 12'h3d0;
		sinewave[432] = 12'h3c4;
		sinewave[433] = 12'h3b9;
		sinewave[434] = 12'h3ae;
		sinewave[435] = 12'h3a3;
		sinewave[436] = 12'h398;
		sinewave[437] = 12'h38d;
		sinewave[438] = 12'h381;
		sinewave[439] = 12'h376;
		sinewave[440] = 12'h36b;
		sinewave[441] = 12'h35f;
		sinewave[442] = 12'h354;
		sinewave[443] = 12'h348;
		sinewave[444] = 12'h33d;
		sinewave[445] = 12'h332;
		sinewave[446] = 12'h326;
		sinewave[447] = 12'h31a;
		sinewave[448] = 12'h30f;
		sinewave[449] = 12'h303;
		sinewave[450] = 12'h2f8;
		sinewave[451] = 12'h2ec;
		sinewave[452] = 12'h2e0;
		sinewave[453] = 12'h2d4;
		sinewave[454] = 12'h2c9;
		sinewave[455] = 12'h2bd;
		sinewave[456] = 12'h2b1;
		sinewave[457] = 12'h2a5;
		sinewave[458] = 12'h299;
		sinewave[459] = 12'h28e;
		sinewave[460] = 12'h282;
		sinewave[461] = 12'h276;
		sinewave[462] = 12'h26a;
		sinewave[463] = 12'h25e;
		sinewave[464] = 12'h252;
		sinewave[465] = 12'h246;
		sinewave[466] = 12'h23a;
		sinewave[467] = 12'h22e;
		sinewave[468] = 12'h221;
		sinewave[469] = 12'h215;
		sinewave[470] = 12'h209;
		sinewave[471] = 12'h1fd;
		sinewave[472] = 12'h1f1;
		sinewave[473] = 12'h1e5;
		sinewave[474] = 12'h1d8;
		sinewave[475] = 12'h1cc;
		sinewave[476] = 12'h1c0;
		sinewave[477] = 12'h1b4;
		sinewave[478] = 12'h1a7;
		sinewave[479] = 12'h19b;
		sinewave[480] = 12'h18f;
		sinewave[481] = 12'h183;
		sinewave[482] = 12'h176;
		sinewave[483] = 12'h16a;
		sinewave[484] = 12'h15d;
		sinewave[485] = 12'h151;
		sinewave[486] = 12'h145;
		sinewave[487] = 12'h138;
		sinewave[488] = 12'h12c;
		sinewave[489] = 12'h11f;
		sinewave[490] = 12'h113;
		sinewave[491] = 12'h107;
		sinewave[492] = 12'hfa;
		sinewave[493] = 12'hee;
		sinewave[494] = 12'he1;
		sinewave[495] = 12'hd5;
		sinewave[496] = 12'hc8;
		sinewave[497] = 12'hbc;
		sinewave[498] = 12'haf;
		sinewave[499] = 12'ha3;
		sinewave[500] = 12'h96;
		sinewave[501] = 12'h8a;
		sinewave[502] = 12'h7d;
		sinewave[503] = 12'h70;
		sinewave[504] = 12'h64;
		sinewave[505] = 12'h57;
		sinewave[506] = 12'h4b;
		sinewave[507] = 12'h3e;
		sinewave[508] = 12'h32;
		sinewave[509] = 12'h25;
		sinewave[510] = 12'h19;
		sinewave[511] = 12'h0c;
		sinewave[512] = 12'h00;
		sinewave[513] = 12'hff4;
		sinewave[514] = 12'hfe7;
		sinewave[515] = 12'hfdb;
		sinewave[516] = 12'hfce;
		sinewave[517] = 12'hfc2;
		sinewave[518] = 12'hfb5;
		sinewave[519] = 12'hfa9;
		sinewave[520] = 12'hf9c;
		sinewave[521] = 12'hf90;
		sinewave[522] = 12'hf83;
		sinewave[523] = 12'hf76;
		sinewave[524] = 12'hf6a;
		sinewave[525] = 12'hf5d;
		sinewave[526] = 12'hf51;
		sinewave[527] = 12'hf44;
		sinewave[528] = 12'hf38;
		sinewave[529] = 12'hf2b;
		sinewave[530] = 12'hf1f;
		sinewave[531] = 12'hf12;
		sinewave[532] = 12'hf06;
		sinewave[533] = 12'hef9;
		sinewave[534] = 12'heed;
		sinewave[535] = 12'hee1;
		sinewave[536] = 12'hed4;
		sinewave[537] = 12'hec8;
		sinewave[538] = 12'hebb;
		sinewave[539] = 12'heaf;
		sinewave[540] = 12'hea3;
		sinewave[541] = 12'he96;
		sinewave[542] = 12'he8a;
		sinewave[543] = 12'he7d;
		sinewave[544] = 12'he71;
		sinewave[545] = 12'he65;
		sinewave[546] = 12'he59;
		sinewave[547] = 12'he4c;
		sinewave[548] = 12'he40;
		sinewave[549] = 12'he34;
		sinewave[550] = 12'he28;
		sinewave[551] = 12'he1b;
		sinewave[552] = 12'he0f;
		sinewave[553] = 12'he03;
		sinewave[554] = 12'hdf7;
		sinewave[555] = 12'hdeb;
		sinewave[556] = 12'hddf;
		sinewave[557] = 12'hdd2;
		sinewave[558] = 12'hdc6;
		sinewave[559] = 12'hdba;
		sinewave[560] = 12'hdae;
		sinewave[561] = 12'hda2;
		sinewave[562] = 12'hd96;
		sinewave[563] = 12'hd8a;
		sinewave[564] = 12'hd7e;
		sinewave[565] = 12'hd72;
		sinewave[566] = 12'hd67;
		sinewave[567] = 12'hd5b;
		sinewave[568] = 12'hd4f;
		sinewave[569] = 12'hd43;
		sinewave[570] = 12'hd37;
		sinewave[571] = 12'hd2c;
		sinewave[572] = 12'hd20;
		sinewave[573] = 12'hd14;
		sinewave[574] = 12'hd08;
		sinewave[575] = 12'hcfd;
		sinewave[576] = 12'hcf1;
		sinewave[577] = 12'hce6;
		sinewave[578] = 12'hcda;
		sinewave[579] = 12'hcce;
		sinewave[580] = 12'hcc3;
		sinewave[581] = 12'hcb8;
		sinewave[582] = 12'hcac;
		sinewave[583] = 12'hca1;
		sinewave[584] = 12'hc95;
		sinewave[585] = 12'hc8a;
		sinewave[586] = 12'hc7f;
		sinewave[587] = 12'hc73;
		sinewave[588] = 12'hc68;
		sinewave[589] = 12'hc5d;
		sinewave[590] = 12'hc52;
		sinewave[591] = 12'hc47;
		sinewave[592] = 12'hc3c;
		sinewave[593] = 12'hc30;
		sinewave[594] = 12'hc25;
		sinewave[595] = 12'hc1a;
		sinewave[596] = 12'hc10;
		sinewave[597] = 12'hc05;
		sinewave[598] = 12'hbfa;
		sinewave[599] = 12'hbef;
		sinewave[600] = 12'hbe4;
		sinewave[601] = 12'hbd9;
		sinewave[602] = 12'hbcf;
		sinewave[603] = 12'hbc4;
		sinewave[604] = 12'hbb9;
		sinewave[605] = 12'hbaf;
		sinewave[606] = 12'hba4;
		sinewave[607] = 12'hb9a;
		sinewave[608] = 12'hb8f;
		sinewave[609] = 12'hb85;
		sinewave[610] = 12'hb7a;
		sinewave[611] = 12'hb70;
		sinewave[612] = 12'hb66;
		sinewave[613] = 12'hb5c;
		sinewave[614] = 12'hb51;
		sinewave[615] = 12'hb47;
		sinewave[616] = 12'hb3d;
		sinewave[617] = 12'hb33;
		sinewave[618] = 12'hb29;
		sinewave[619] = 12'hb1f;
		sinewave[620] = 12'hb15;
		sinewave[621] = 12'hb0b;
		sinewave[622] = 12'hb01;
		sinewave[623] = 12'haf8;
		sinewave[624] = 12'haee;
		sinewave[625] = 12'hae4;
		sinewave[626] = 12'hadb;
		sinewave[627] = 12'had1;
		sinewave[628] = 12'hac7;
		sinewave[629] = 12'habe;
		sinewave[630] = 12'hab5;
		sinewave[631] = 12'haab;
		sinewave[632] = 12'haa2;
		sinewave[633] = 12'ha99;
		sinewave[634] = 12'ha8f;
		sinewave[635] = 12'ha86;
		sinewave[636] = 12'ha7d;
		sinewave[637] = 12'ha74;
		sinewave[638] = 12'ha6b;
		sinewave[639] = 12'ha62;
		sinewave[640] = 12'ha59;
		sinewave[641] = 12'ha50;
		sinewave[642] = 12'ha47;
		sinewave[643] = 12'ha3f;
		sinewave[644] = 12'ha36;
		sinewave[645] = 12'ha2d;
		sinewave[646] = 12'ha25;
		sinewave[647] = 12'ha1c;
		sinewave[648] = 12'ha14;
		sinewave[649] = 12'ha0b;
		sinewave[650] = 12'ha03;
		sinewave[651] = 12'h9fb;
		sinewave[652] = 12'h9f2;
		sinewave[653] = 12'h9ea;
		sinewave[654] = 12'h9e2;
		sinewave[655] = 12'h9da;
		sinewave[656] = 12'h9d2;
		sinewave[657] = 12'h9ca;
		sinewave[658] = 12'h9c2;
		sinewave[659] = 12'h9bb;
		sinewave[660] = 12'h9b3;
		sinewave[661] = 12'h9ab;
		sinewave[662] = 12'h9a3;
		sinewave[663] = 12'h99c;
		sinewave[664] = 12'h994;
		sinewave[665] = 12'h98d;
		sinewave[666] = 12'h985;
		sinewave[667] = 12'h97e;
		sinewave[668] = 12'h977;
		sinewave[669] = 12'h970;
		sinewave[670] = 12'h969;
		sinewave[671] = 12'h961;
		sinewave[672] = 12'h95a;
		sinewave[673] = 12'h954;
		sinewave[674] = 12'h94d;
		sinewave[675] = 12'h946;
		sinewave[676] = 12'h93f;
		sinewave[677] = 12'h938;
		sinewave[678] = 12'h932;
		sinewave[679] = 12'h92b;
		sinewave[680] = 12'h925;
		sinewave[681] = 12'h91e;
		sinewave[682] = 12'h918;
		sinewave[683] = 12'h912;
		sinewave[684] = 12'h90b;
		sinewave[685] = 12'h905;
		sinewave[686] = 12'h8ff;
		sinewave[687] = 12'h8f9;
		sinewave[688] = 12'h8f3;
		sinewave[689] = 12'h8ed;
		sinewave[690] = 12'h8e8;
		sinewave[691] = 12'h8e2;
		sinewave[692] = 12'h8dc;
		sinewave[693] = 12'h8d6;
		sinewave[694] = 12'h8d1;
		sinewave[695] = 12'h8cb;
		sinewave[696] = 12'h8c6;
		sinewave[697] = 12'h8c1;
		sinewave[698] = 12'h8bb;
		sinewave[699] = 12'h8b6;
		sinewave[700] = 12'h8b1;
		sinewave[701] = 12'h8ac;
		sinewave[702] = 12'h8a7;
		sinewave[703] = 12'h8a2;
		sinewave[704] = 12'h89d;
		sinewave[705] = 12'h899;
		sinewave[706] = 12'h894;
		sinewave[707] = 12'h88f;
		sinewave[708] = 12'h88b;
		sinewave[709] = 12'h886;
		sinewave[710] = 12'h882;
		sinewave[711] = 12'h87d;
		sinewave[712] = 12'h879;
		sinewave[713] = 12'h875;
		sinewave[714] = 12'h871;
		sinewave[715] = 12'h86d;
		sinewave[716] = 12'h869;
		sinewave[717] = 12'h865;
		sinewave[718] = 12'h861;
		sinewave[719] = 12'h85d;
		sinewave[720] = 12'h85a;
		sinewave[721] = 12'h856;
		sinewave[722] = 12'h852;
		sinewave[723] = 12'h84f;
		sinewave[724] = 12'h84c;
		sinewave[725] = 12'h848;
		sinewave[726] = 12'h845;
		sinewave[727] = 12'h842;
		sinewave[728] = 12'h83f;
		sinewave[729] = 12'h83c;
		sinewave[730] = 12'h839;
		sinewave[731] = 12'h836;
		sinewave[732] = 12'h833;
		sinewave[733] = 12'h831;
		sinewave[734] = 12'h82e;
		sinewave[735] = 12'h82b;
		sinewave[736] = 12'h829;
		sinewave[737] = 12'h826;
		sinewave[738] = 12'h824;
		sinewave[739] = 12'h822;
		sinewave[740] = 12'h820;
		sinewave[741] = 12'h81e;
		sinewave[742] = 12'h81b;
		sinewave[743] = 12'h81a;
		sinewave[744] = 12'h818;
		sinewave[745] = 12'h816;
		sinewave[746] = 12'h814;
		sinewave[747] = 12'h812;
		sinewave[748] = 12'h811;
		sinewave[749] = 12'h80f;
		sinewave[750] = 12'h80e;
		sinewave[751] = 12'h80d;
		sinewave[752] = 12'h80b;
		sinewave[753] = 12'h80a;
		sinewave[754] = 12'h809;
		sinewave[755] = 12'h808;
		sinewave[756] = 12'h807;
		sinewave[757] = 12'h806;
		sinewave[758] = 12'h805;
		sinewave[759] = 12'h805;
		sinewave[760] = 12'h804;
		sinewave[761] = 12'h803;
		sinewave[762] = 12'h803;
		sinewave[763] = 12'h802;
		sinewave[764] = 12'h802;
		sinewave[765] = 12'h802;
		sinewave[766] = 12'h802;
		sinewave[767] = 12'h802;
		sinewave[768] = 12'h801;
		sinewave[769] = 12'h802;
		sinewave[770] = 12'h802;
		sinewave[771] = 12'h802;
		sinewave[772] = 12'h802;
		sinewave[773] = 12'h802;
		sinewave[774] = 12'h803;
		sinewave[775] = 12'h803;
		sinewave[776] = 12'h804;
		sinewave[777] = 12'h805;
		sinewave[778] = 12'h805;
		sinewave[779] = 12'h806;
		sinewave[780] = 12'h807;
		sinewave[781] = 12'h808;
		sinewave[782] = 12'h809;
		sinewave[783] = 12'h80a;
		sinewave[784] = 12'h80b;
		sinewave[785] = 12'h80d;
		sinewave[786] = 12'h80e;
		sinewave[787] = 12'h80f;
		sinewave[788] = 12'h811;
		sinewave[789] = 12'h812;
		sinewave[790] = 12'h814;
		sinewave[791] = 12'h816;
		sinewave[792] = 12'h818;
		sinewave[793] = 12'h81a;
		sinewave[794] = 12'h81b;
		sinewave[795] = 12'h81e;
		sinewave[796] = 12'h820;
		sinewave[797] = 12'h822;
		sinewave[798] = 12'h824;
		sinewave[799] = 12'h826;
		sinewave[800] = 12'h829;
		sinewave[801] = 12'h82b;
		sinewave[802] = 12'h82e;
		sinewave[803] = 12'h831;
		sinewave[804] = 12'h833;
		sinewave[805] = 12'h836;
		sinewave[806] = 12'h839;
		sinewave[807] = 12'h83c;
		sinewave[808] = 12'h83f;
		sinewave[809] = 12'h842;
		sinewave[810] = 12'h845;
		sinewave[811] = 12'h848;
		sinewave[812] = 12'h84c;
		sinewave[813] = 12'h84f;
		sinewave[814] = 12'h852;
		sinewave[815] = 12'h856;
		sinewave[816] = 12'h85a;
		sinewave[817] = 12'h85d;
		sinewave[818] = 12'h861;
		sinewave[819] = 12'h865;
		sinewave[820] = 12'h869;
		sinewave[821] = 12'h86d;
		sinewave[822] = 12'h871;
		sinewave[823] = 12'h875;
		sinewave[824] = 12'h879;
		sinewave[825] = 12'h87d;
		sinewave[826] = 12'h882;
		sinewave[827] = 12'h886;
		sinewave[828] = 12'h88b;
		sinewave[829] = 12'h88f;
		sinewave[830] = 12'h894;
		sinewave[831] = 12'h899;
		sinewave[832] = 12'h89d;
		sinewave[833] = 12'h8a2;
		sinewave[834] = 12'h8a7;
		sinewave[835] = 12'h8ac;
		sinewave[836] = 12'h8b1;
		sinewave[837] = 12'h8b6;
		sinewave[838] = 12'h8bb;
		sinewave[839] = 12'h8c1;
		sinewave[840] = 12'h8c6;
		sinewave[841] = 12'h8cb;
		sinewave[842] = 12'h8d1;
		sinewave[843] = 12'h8d6;
		sinewave[844] = 12'h8dc;
		sinewave[845] = 12'h8e2;
		sinewave[846] = 12'h8e8;
		sinewave[847] = 12'h8ed;
		sinewave[848] = 12'h8f3;
		sinewave[849] = 12'h8f9;
		sinewave[850] = 12'h8ff;
		sinewave[851] = 12'h905;
		sinewave[852] = 12'h90b;
		sinewave[853] = 12'h912;
		sinewave[854] = 12'h918;
		sinewave[855] = 12'h91e;
		sinewave[856] = 12'h925;
		sinewave[857] = 12'h92b;
		sinewave[858] = 12'h932;
		sinewave[859] = 12'h938;
		sinewave[860] = 12'h93f;
		sinewave[861] = 12'h946;
		sinewave[862] = 12'h94d;
		sinewave[863] = 12'h954;
		sinewave[864] = 12'h95a;
		sinewave[865] = 12'h961;
		sinewave[866] = 12'h969;
		sinewave[867] = 12'h970;
		sinewave[868] = 12'h977;
		sinewave[869] = 12'h97e;
		sinewave[870] = 12'h985;
		sinewave[871] = 12'h98d;
		sinewave[872] = 12'h994;
		sinewave[873] = 12'h99c;
		sinewave[874] = 12'h9a3;
		sinewave[875] = 12'h9ab;
		sinewave[876] = 12'h9b3;
		sinewave[877] = 12'h9bb;
		sinewave[878] = 12'h9c2;
		sinewave[879] = 12'h9ca;
		sinewave[880] = 12'h9d2;
		sinewave[881] = 12'h9da;
		sinewave[882] = 12'h9e2;
		sinewave[883] = 12'h9ea;
		sinewave[884] = 12'h9f2;
		sinewave[885] = 12'h9fb;
		sinewave[886] = 12'ha03;
		sinewave[887] = 12'ha0b;
		sinewave[888] = 12'ha14;
		sinewave[889] = 12'ha1c;
		sinewave[890] = 12'ha25;
		sinewave[891] = 12'ha2d;
		sinewave[892] = 12'ha36;
		sinewave[893] = 12'ha3f;
		sinewave[894] = 12'ha47;
		sinewave[895] = 12'ha50;
		sinewave[896] = 12'ha59;
		sinewave[897] = 12'ha62;
		sinewave[898] = 12'ha6b;
		sinewave[899] = 12'ha74;
		sinewave[900] = 12'ha7d;
		sinewave[901] = 12'ha86;
		sinewave[902] = 12'ha8f;
		sinewave[903] = 12'ha99;
		sinewave[904] = 12'haa2;
		sinewave[905] = 12'haab;
		sinewave[906] = 12'hab5;
		sinewave[907] = 12'habe;
		sinewave[908] = 12'hac7;
		sinewave[909] = 12'had1;
		sinewave[910] = 12'hadb;
		sinewave[911] = 12'hae4;
		sinewave[912] = 12'haee;
		sinewave[913] = 12'haf8;
		sinewave[914] = 12'hb01;
		sinewave[915] = 12'hb0b;
		sinewave[916] = 12'hb15;
		sinewave[917] = 12'hb1f;
		sinewave[918] = 12'hb29;
		sinewave[919] = 12'hb33;
		sinewave[920] = 12'hb3d;
		sinewave[921] = 12'hb47;
		sinewave[922] = 12'hb51;
		sinewave[923] = 12'hb5c;
		sinewave[924] = 12'hb66;
		sinewave[925] = 12'hb70;
		sinewave[926] = 12'hb7a;
		sinewave[927] = 12'hb85;
		sinewave[928] = 12'hb8f;
		sinewave[929] = 12'hb9a;
		sinewave[930] = 12'hba4;
		sinewave[931] = 12'hbaf;
		sinewave[932] = 12'hbb9;
		sinewave[933] = 12'hbc4;
		sinewave[934] = 12'hbcf;
		sinewave[935] = 12'hbd9;
		sinewave[936] = 12'hbe4;
		sinewave[937] = 12'hbef;
		sinewave[938] = 12'hbfa;
		sinewave[939] = 12'hc05;
		sinewave[940] = 12'hc10;
		sinewave[941] = 12'hc1a;
		sinewave[942] = 12'hc25;
		sinewave[943] = 12'hc30;
		sinewave[944] = 12'hc3c;
		sinewave[945] = 12'hc47;
		sinewave[946] = 12'hc52;
		sinewave[947] = 12'hc5d;
		sinewave[948] = 12'hc68;
		sinewave[949] = 12'hc73;
		sinewave[950] = 12'hc7f;
		sinewave[951] = 12'hc8a;
		sinewave[952] = 12'hc95;
		sinewave[953] = 12'hca1;
		sinewave[954] = 12'hcac;
		sinewave[955] = 12'hcb8;
		sinewave[956] = 12'hcc3;
		sinewave[957] = 12'hcce;
		sinewave[958] = 12'hcda;
		sinewave[959] = 12'hce6;
		sinewave[960] = 12'hcf1;
		sinewave[961] = 12'hcfd;
		sinewave[962] = 12'hd08;
		sinewave[963] = 12'hd14;
		sinewave[964] = 12'hd20;
		sinewave[965] = 12'hd2c;
		sinewave[966] = 12'hd37;
		sinewave[967] = 12'hd43;
		sinewave[968] = 12'hd4f;
		sinewave[969] = 12'hd5b;
		sinewave[970] = 12'hd67;
		sinewave[971] = 12'hd72;
		sinewave[972] = 12'hd7e;
		sinewave[973] = 12'hd8a;
		sinewave[974] = 12'hd96;
		sinewave[975] = 12'hda2;
		sinewave[976] = 12'hdae;
		sinewave[977] = 12'hdba;
		sinewave[978] = 12'hdc6;
		sinewave[979] = 12'hdd2;
		sinewave[980] = 12'hddf;
		sinewave[981] = 12'hdeb;
		sinewave[982] = 12'hdf7;
		sinewave[983] = 12'he03;
		sinewave[984] = 12'he0f;
		sinewave[985] = 12'he1b;
		sinewave[986] = 12'he28;
		sinewave[987] = 12'he34;
		sinewave[988] = 12'he40;
		sinewave[989] = 12'he4c;
		sinewave[990] = 12'he59;
		sinewave[991] = 12'he65;
		sinewave[992] = 12'he71;
		sinewave[993] = 12'he7d;
		sinewave[994] = 12'he8a;
		sinewave[995] = 12'he96;
		sinewave[996] = 12'hea3;
		sinewave[997] = 12'heaf;
		sinewave[998] = 12'hebb;
		sinewave[999] = 12'hec8;
		sinewave[1000] = 12'hed4;
		sinewave[1001] = 12'hee1;
		sinewave[1002] = 12'heed;
		sinewave[1003] = 12'hef9;
		sinewave[1004] = 12'hf06;
		sinewave[1005] = 12'hf12;
		sinewave[1006] = 12'hf1f;
		sinewave[1007] = 12'hf2b;
		sinewave[1008] = 12'hf38;
		sinewave[1009] = 12'hf44;
		sinewave[1010] = 12'hf51;
		sinewave[1011] = 12'hf5d;
		sinewave[1012] = 12'hf6a;
		sinewave[1013] = 12'hf76;
		sinewave[1014] = 12'hf83;
		sinewave[1015] = 12'hf90;
		sinewave[1016] = 12'hf9c;
		sinewave[1017] = 12'hfa9;
		sinewave[1018] = 12'hfb5;
		sinewave[1019] = 12'hfc2;
		sinewave[1020] = 12'hfce;
		sinewave[1021] = 12'hfdb;
		sinewave[1022] = 12'hfe7;
		sinewave[1023] = 12'hff4;
	end
	
	// === SAMPLER ===
	always @(posedge inCLK) begin
		// Perform phase update and sample output shift only when sampling is clock-enabled
		if (inSampleClockCE) begin
			phase <= phase + frequency_step[inMidiFrequencyIndex];
			
			// Switch on sample wave mode
			case(inWaveMode)
				// 0 - Sinewave: signed 12 bit Sinewave lookup table from 10 phase bits (1024 unique sinewave samples)
				0: outSample <= sinewave[phase[N-1:N-10]];
				// 1 - Squarewave: signed 12 bit positive and negative maximums
				1: outSample <= (phase[N-1] ?  12'h801 : 12'h7ff); 
				// default - Sinewave
				default: outSample <= sinewave[phase[N-1:N-10]];
			endcase
		end
	end
endmodule
