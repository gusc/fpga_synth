`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:56:17 06/14/2018 
// Design Name: 
// Module Name:    tableSinewave 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module tableSinewave(idx, sinewave);
input [9:0] idx;
output reg [11:0] sinewave = 0;
always @(idx) begin

	// Samples: 1024
	// Top value: 2047
	// Mid value: 0
	// Bottom value: -2047
	case(idx)
	10'd0   : sinewave = 12'h00;
	10'd1   : sinewave = 12'h0c;
	10'd2   : sinewave = 12'h19;
	10'd3   : sinewave = 12'h25;
	10'd4   : sinewave = 12'h32;
	10'd5   : sinewave = 12'h3e;
	10'd6   : sinewave = 12'h4b;
	10'd7   : sinewave = 12'h57;
	10'd8   : sinewave = 12'h64;
	10'd9   : sinewave = 12'h70;
	10'd10  : sinewave = 12'h7d;
	10'd11  : sinewave = 12'h8a;
	10'd12  : sinewave = 12'h96;
	10'd13  : sinewave = 12'ha3;
	10'd14  : sinewave = 12'haf;
	10'd15  : sinewave = 12'hbc;
	10'd16  : sinewave = 12'hc8;
	10'd17  : sinewave = 12'hd5;
	10'd18  : sinewave = 12'he1;
	10'd19  : sinewave = 12'hee;
	10'd20  : sinewave = 12'hfa;
	10'd21  : sinewave = 12'h107;
	10'd22  : sinewave = 12'h113;
	10'd23  : sinewave = 12'h11f;
	10'd24  : sinewave = 12'h12c;
	10'd25  : sinewave = 12'h138;
	10'd26  : sinewave = 12'h145;
	10'd27  : sinewave = 12'h151;
	10'd28  : sinewave = 12'h15d;
	10'd29  : sinewave = 12'h16a;
	10'd30  : sinewave = 12'h176;
	10'd31  : sinewave = 12'h183;
	10'd32  : sinewave = 12'h18f;
	10'd33  : sinewave = 12'h19b;
	10'd34  : sinewave = 12'h1a7;
	10'd35  : sinewave = 12'h1b4;
	10'd36  : sinewave = 12'h1c0;
	10'd37  : sinewave = 12'h1cc;
	10'd38  : sinewave = 12'h1d8;
	10'd39  : sinewave = 12'h1e5;
	10'd40  : sinewave = 12'h1f1;
	10'd41  : sinewave = 12'h1fd;
	10'd42  : sinewave = 12'h209;
	10'd43  : sinewave = 12'h215;
	10'd44  : sinewave = 12'h221;
	10'd45  : sinewave = 12'h22e;
	10'd46  : sinewave = 12'h23a;
	10'd47  : sinewave = 12'h246;
	10'd48  : sinewave = 12'h252;
	10'd49  : sinewave = 12'h25e;
	10'd50  : sinewave = 12'h26a;
	10'd51  : sinewave = 12'h276;
	10'd52  : sinewave = 12'h282;
	10'd53  : sinewave = 12'h28e;
	10'd54  : sinewave = 12'h299;
	10'd55  : sinewave = 12'h2a5;
	10'd56  : sinewave = 12'h2b1;
	10'd57  : sinewave = 12'h2bd;
	10'd58  : sinewave = 12'h2c9;
	10'd59  : sinewave = 12'h2d4;
	10'd60  : sinewave = 12'h2e0;
	10'd61  : sinewave = 12'h2ec;
	10'd62  : sinewave = 12'h2f8;
	10'd63  : sinewave = 12'h303;
	10'd64  : sinewave = 12'h30f;
	10'd65  : sinewave = 12'h31a;
	10'd66  : sinewave = 12'h326;
	10'd67  : sinewave = 12'h332;
	10'd68  : sinewave = 12'h33d;
	10'd69  : sinewave = 12'h348;
	10'd70  : sinewave = 12'h354;
	10'd71  : sinewave = 12'h35f;
	10'd72  : sinewave = 12'h36b;
	10'd73  : sinewave = 12'h376;
	10'd74  : sinewave = 12'h381;
	10'd75  : sinewave = 12'h38d;
	10'd76  : sinewave = 12'h398;
	10'd77  : sinewave = 12'h3a3;
	10'd78  : sinewave = 12'h3ae;
	10'd79  : sinewave = 12'h3b9;
	10'd80  : sinewave = 12'h3c4;
	10'd81  : sinewave = 12'h3d0;
	10'd82  : sinewave = 12'h3db;
	10'd83  : sinewave = 12'h3e6;
	10'd84  : sinewave = 12'h3f0;
	10'd85  : sinewave = 12'h3fb;
	10'd86  : sinewave = 12'h406;
	10'd87  : sinewave = 12'h411;
	10'd88  : sinewave = 12'h41c;
	10'd89  : sinewave = 12'h427;
	10'd90  : sinewave = 12'h431;
	10'd91  : sinewave = 12'h43c;
	10'd92  : sinewave = 12'h447;
	10'd93  : sinewave = 12'h451;
	10'd94  : sinewave = 12'h45c;
	10'd95  : sinewave = 12'h466;
	10'd96  : sinewave = 12'h471;
	10'd97  : sinewave = 12'h47b;
	10'd98  : sinewave = 12'h486;
	10'd99  : sinewave = 12'h490;
	10'd100 : sinewave = 12'h49a;
	10'd101 : sinewave = 12'h4a4;
	10'd102 : sinewave = 12'h4af;
	10'd103 : sinewave = 12'h4b9;
	10'd104 : sinewave = 12'h4c3;
	10'd105 : sinewave = 12'h4cd;
	10'd106 : sinewave = 12'h4d7;
	10'd107 : sinewave = 12'h4e1;
	10'd108 : sinewave = 12'h4eb;
	10'd109 : sinewave = 12'h4f5;
	10'd110 : sinewave = 12'h4ff;
	10'd111 : sinewave = 12'h508;
	10'd112 : sinewave = 12'h512;
	10'd113 : sinewave = 12'h51c;
	10'd114 : sinewave = 12'h525;
	10'd115 : sinewave = 12'h52f;
	10'd116 : sinewave = 12'h539;
	10'd117 : sinewave = 12'h542;
	10'd118 : sinewave = 12'h54b;
	10'd119 : sinewave = 12'h555;
	10'd120 : sinewave = 12'h55e;
	10'd121 : sinewave = 12'h567;
	10'd122 : sinewave = 12'h571;
	10'd123 : sinewave = 12'h57a;
	10'd124 : sinewave = 12'h583;
	10'd125 : sinewave = 12'h58c;
	10'd126 : sinewave = 12'h595;
	10'd127 : sinewave = 12'h59e;
	10'd128 : sinewave = 12'h5a7;
	10'd129 : sinewave = 12'h5b0;
	10'd130 : sinewave = 12'h5b9;
	10'd131 : sinewave = 12'h5c1;
	10'd132 : sinewave = 12'h5ca;
	10'd133 : sinewave = 12'h5d3;
	10'd134 : sinewave = 12'h5db;
	10'd135 : sinewave = 12'h5e4;
	10'd136 : sinewave = 12'h5ec;
	10'd137 : sinewave = 12'h5f5;
	10'd138 : sinewave = 12'h5fd;
	10'd139 : sinewave = 12'h605;
	10'd140 : sinewave = 12'h60e;
	10'd141 : sinewave = 12'h616;
	10'd142 : sinewave = 12'h61e;
	10'd143 : sinewave = 12'h626;
	10'd144 : sinewave = 12'h62e;
	10'd145 : sinewave = 12'h636;
	10'd146 : sinewave = 12'h63e;
	10'd147 : sinewave = 12'h645;
	10'd148 : sinewave = 12'h64d;
	10'd149 : sinewave = 12'h655;
	10'd150 : sinewave = 12'h65d;
	10'd151 : sinewave = 12'h664;
	10'd152 : sinewave = 12'h66c;
	10'd153 : sinewave = 12'h673;
	10'd154 : sinewave = 12'h67b;
	10'd155 : sinewave = 12'h682;
	10'd156 : sinewave = 12'h689;
	10'd157 : sinewave = 12'h690;
	10'd158 : sinewave = 12'h697;
	10'd159 : sinewave = 12'h69f;
	10'd160 : sinewave = 12'h6a6;
	10'd161 : sinewave = 12'h6ac;
	10'd162 : sinewave = 12'h6b3;
	10'd163 : sinewave = 12'h6ba;
	10'd164 : sinewave = 12'h6c1;
	10'd165 : sinewave = 12'h6c8;
	10'd166 : sinewave = 12'h6ce;
	10'd167 : sinewave = 12'h6d5;
	10'd168 : sinewave = 12'h6db;
	10'd169 : sinewave = 12'h6e2;
	10'd170 : sinewave = 12'h6e8;
	10'd171 : sinewave = 12'h6ee;
	10'd172 : sinewave = 12'h6f5;
	10'd173 : sinewave = 12'h6fb;
	10'd174 : sinewave = 12'h701;
	10'd175 : sinewave = 12'h707;
	10'd176 : sinewave = 12'h70d;
	10'd177 : sinewave = 12'h713;
	10'd178 : sinewave = 12'h718;
	10'd179 : sinewave = 12'h71e;
	10'd180 : sinewave = 12'h724;
	10'd181 : sinewave = 12'h72a;
	10'd182 : sinewave = 12'h72f;
	10'd183 : sinewave = 12'h735;
	10'd184 : sinewave = 12'h73a;
	10'd185 : sinewave = 12'h73f;
	10'd186 : sinewave = 12'h745;
	10'd187 : sinewave = 12'h74a;
	10'd188 : sinewave = 12'h74f;
	10'd189 : sinewave = 12'h754;
	10'd190 : sinewave = 12'h759;
	10'd191 : sinewave = 12'h75e;
	10'd192 : sinewave = 12'h763;
	10'd193 : sinewave = 12'h767;
	10'd194 : sinewave = 12'h76c;
	10'd195 : sinewave = 12'h771;
	10'd196 : sinewave = 12'h775;
	10'd197 : sinewave = 12'h77a;
	10'd198 : sinewave = 12'h77e;
	10'd199 : sinewave = 12'h783;
	10'd200 : sinewave = 12'h787;
	10'd201 : sinewave = 12'h78b;
	10'd202 : sinewave = 12'h78f;
	10'd203 : sinewave = 12'h793;
	10'd204 : sinewave = 12'h797;
	10'd205 : sinewave = 12'h79b;
	10'd206 : sinewave = 12'h79f;
	10'd207 : sinewave = 12'h7a3;
	10'd208 : sinewave = 12'h7a6;
	10'd209 : sinewave = 12'h7aa;
	10'd210 : sinewave = 12'h7ae;
	10'd211 : sinewave = 12'h7b1;
	10'd212 : sinewave = 12'h7b4;
	10'd213 : sinewave = 12'h7b8;
	10'd214 : sinewave = 12'h7bb;
	10'd215 : sinewave = 12'h7be;
	10'd216 : sinewave = 12'h7c1;
	10'd217 : sinewave = 12'h7c4;
	10'd218 : sinewave = 12'h7c7;
	10'd219 : sinewave = 12'h7ca;
	10'd220 : sinewave = 12'h7cd;
	10'd221 : sinewave = 12'h7cf;
	10'd222 : sinewave = 12'h7d2;
	10'd223 : sinewave = 12'h7d5;
	10'd224 : sinewave = 12'h7d7;
	10'd225 : sinewave = 12'h7da;
	10'd226 : sinewave = 12'h7dc;
	10'd227 : sinewave = 12'h7de;
	10'd228 : sinewave = 12'h7e0;
	10'd229 : sinewave = 12'h7e2;
	10'd230 : sinewave = 12'h7e5;
	10'd231 : sinewave = 12'h7e6;
	10'd232 : sinewave = 12'h7e8;
	10'd233 : sinewave = 12'h7ea;
	10'd234 : sinewave = 12'h7ec;
	10'd235 : sinewave = 12'h7ee;
	10'd236 : sinewave = 12'h7ef;
	10'd237 : sinewave = 12'h7f1;
	10'd238 : sinewave = 12'h7f2;
	10'd239 : sinewave = 12'h7f3;
	10'd240 : sinewave = 12'h7f5;
	10'd241 : sinewave = 12'h7f6;
	10'd242 : sinewave = 12'h7f7;
	10'd243 : sinewave = 12'h7f8;
	10'd244 : sinewave = 12'h7f9;
	10'd245 : sinewave = 12'h7fa;
	10'd246 : sinewave = 12'h7fb;
	10'd247 : sinewave = 12'h7fb;
	10'd248 : sinewave = 12'h7fc;
	10'd249 : sinewave = 12'h7fd;
	10'd250 : sinewave = 12'h7fd;
	10'd251 : sinewave = 12'h7fe;
	10'd252 : sinewave = 12'h7fe;
	10'd253 : sinewave = 12'h7fe;
	10'd254 : sinewave = 12'h7fe;
	10'd255 : sinewave = 12'h7fe;
	10'd256 : sinewave = 12'h7ff;
	10'd257 : sinewave = 12'h7fe;
	10'd258 : sinewave = 12'h7fe;
	10'd259 : sinewave = 12'h7fe;
	10'd260 : sinewave = 12'h7fe;
	10'd261 : sinewave = 12'h7fe;
	10'd262 : sinewave = 12'h7fd;
	10'd263 : sinewave = 12'h7fd;
	10'd264 : sinewave = 12'h7fc;
	10'd265 : sinewave = 12'h7fb;
	10'd266 : sinewave = 12'h7fb;
	10'd267 : sinewave = 12'h7fa;
	10'd268 : sinewave = 12'h7f9;
	10'd269 : sinewave = 12'h7f8;
	10'd270 : sinewave = 12'h7f7;
	10'd271 : sinewave = 12'h7f6;
	10'd272 : sinewave = 12'h7f5;
	10'd273 : sinewave = 12'h7f3;
	10'd274 : sinewave = 12'h7f2;
	10'd275 : sinewave = 12'h7f1;
	10'd276 : sinewave = 12'h7ef;
	10'd277 : sinewave = 12'h7ee;
	10'd278 : sinewave = 12'h7ec;
	10'd279 : sinewave = 12'h7ea;
	10'd280 : sinewave = 12'h7e8;
	10'd281 : sinewave = 12'h7e6;
	10'd282 : sinewave = 12'h7e5;
	10'd283 : sinewave = 12'h7e2;
	10'd284 : sinewave = 12'h7e0;
	10'd285 : sinewave = 12'h7de;
	10'd286 : sinewave = 12'h7dc;
	10'd287 : sinewave = 12'h7da;
	10'd288 : sinewave = 12'h7d7;
	10'd289 : sinewave = 12'h7d5;
	10'd290 : sinewave = 12'h7d2;
	10'd291 : sinewave = 12'h7cf;
	10'd292 : sinewave = 12'h7cd;
	10'd293 : sinewave = 12'h7ca;
	10'd294 : sinewave = 12'h7c7;
	10'd295 : sinewave = 12'h7c4;
	10'd296 : sinewave = 12'h7c1;
	10'd297 : sinewave = 12'h7be;
	10'd298 : sinewave = 12'h7bb;
	10'd299 : sinewave = 12'h7b8;
	10'd300 : sinewave = 12'h7b4;
	10'd301 : sinewave = 12'h7b1;
	10'd302 : sinewave = 12'h7ae;
	10'd303 : sinewave = 12'h7aa;
	10'd304 : sinewave = 12'h7a6;
	10'd305 : sinewave = 12'h7a3;
	10'd306 : sinewave = 12'h79f;
	10'd307 : sinewave = 12'h79b;
	10'd308 : sinewave = 12'h797;
	10'd309 : sinewave = 12'h793;
	10'd310 : sinewave = 12'h78f;
	10'd311 : sinewave = 12'h78b;
	10'd312 : sinewave = 12'h787;
	10'd313 : sinewave = 12'h783;
	10'd314 : sinewave = 12'h77e;
	10'd315 : sinewave = 12'h77a;
	10'd316 : sinewave = 12'h775;
	10'd317 : sinewave = 12'h771;
	10'd318 : sinewave = 12'h76c;
	10'd319 : sinewave = 12'h767;
	10'd320 : sinewave = 12'h763;
	10'd321 : sinewave = 12'h75e;
	10'd322 : sinewave = 12'h759;
	10'd323 : sinewave = 12'h754;
	10'd324 : sinewave = 12'h74f;
	10'd325 : sinewave = 12'h74a;
	10'd326 : sinewave = 12'h745;
	10'd327 : sinewave = 12'h73f;
	10'd328 : sinewave = 12'h73a;
	10'd329 : sinewave = 12'h735;
	10'd330 : sinewave = 12'h72f;
	10'd331 : sinewave = 12'h72a;
	10'd332 : sinewave = 12'h724;
	10'd333 : sinewave = 12'h71e;
	10'd334 : sinewave = 12'h718;
	10'd335 : sinewave = 12'h713;
	10'd336 : sinewave = 12'h70d;
	10'd337 : sinewave = 12'h707;
	10'd338 : sinewave = 12'h701;
	10'd339 : sinewave = 12'h6fb;
	10'd340 : sinewave = 12'h6f5;
	10'd341 : sinewave = 12'h6ee;
	10'd342 : sinewave = 12'h6e8;
	10'd343 : sinewave = 12'h6e2;
	10'd344 : sinewave = 12'h6db;
	10'd345 : sinewave = 12'h6d5;
	10'd346 : sinewave = 12'h6ce;
	10'd347 : sinewave = 12'h6c8;
	10'd348 : sinewave = 12'h6c1;
	10'd349 : sinewave = 12'h6ba;
	10'd350 : sinewave = 12'h6b3;
	10'd351 : sinewave = 12'h6ac;
	10'd352 : sinewave = 12'h6a6;
	10'd353 : sinewave = 12'h69f;
	10'd354 : sinewave = 12'h697;
	10'd355 : sinewave = 12'h690;
	10'd356 : sinewave = 12'h689;
	10'd357 : sinewave = 12'h682;
	10'd358 : sinewave = 12'h67b;
	10'd359 : sinewave = 12'h673;
	10'd360 : sinewave = 12'h66c;
	10'd361 : sinewave = 12'h664;
	10'd362 : sinewave = 12'h65d;
	10'd363 : sinewave = 12'h655;
	10'd364 : sinewave = 12'h64d;
	10'd365 : sinewave = 12'h645;
	10'd366 : sinewave = 12'h63e;
	10'd367 : sinewave = 12'h636;
	10'd368 : sinewave = 12'h62e;
	10'd369 : sinewave = 12'h626;
	10'd370 : sinewave = 12'h61e;
	10'd371 : sinewave = 12'h616;
	10'd372 : sinewave = 12'h60e;
	10'd373 : sinewave = 12'h605;
	10'd374 : sinewave = 12'h5fd;
	10'd375 : sinewave = 12'h5f5;
	10'd376 : sinewave = 12'h5ec;
	10'd377 : sinewave = 12'h5e4;
	10'd378 : sinewave = 12'h5db;
	10'd379 : sinewave = 12'h5d3;
	10'd380 : sinewave = 12'h5ca;
	10'd381 : sinewave = 12'h5c1;
	10'd382 : sinewave = 12'h5b9;
	10'd383 : sinewave = 12'h5b0;
	10'd384 : sinewave = 12'h5a7;
	10'd385 : sinewave = 12'h59e;
	10'd386 : sinewave = 12'h595;
	10'd387 : sinewave = 12'h58c;
	10'd388 : sinewave = 12'h583;
	10'd389 : sinewave = 12'h57a;
	10'd390 : sinewave = 12'h571;
	10'd391 : sinewave = 12'h567;
	10'd392 : sinewave = 12'h55e;
	10'd393 : sinewave = 12'h555;
	10'd394 : sinewave = 12'h54b;
	10'd395 : sinewave = 12'h542;
	10'd396 : sinewave = 12'h539;
	10'd397 : sinewave = 12'h52f;
	10'd398 : sinewave = 12'h525;
	10'd399 : sinewave = 12'h51c;
	10'd400 : sinewave = 12'h512;
	10'd401 : sinewave = 12'h508;
	10'd402 : sinewave = 12'h4ff;
	10'd403 : sinewave = 12'h4f5;
	10'd404 : sinewave = 12'h4eb;
	10'd405 : sinewave = 12'h4e1;
	10'd406 : sinewave = 12'h4d7;
	10'd407 : sinewave = 12'h4cd;
	10'd408 : sinewave = 12'h4c3;
	10'd409 : sinewave = 12'h4b9;
	10'd410 : sinewave = 12'h4af;
	10'd411 : sinewave = 12'h4a4;
	10'd412 : sinewave = 12'h49a;
	10'd413 : sinewave = 12'h490;
	10'd414 : sinewave = 12'h486;
	10'd415 : sinewave = 12'h47b;
	10'd416 : sinewave = 12'h471;
	10'd417 : sinewave = 12'h466;
	10'd418 : sinewave = 12'h45c;
	10'd419 : sinewave = 12'h451;
	10'd420 : sinewave = 12'h447;
	10'd421 : sinewave = 12'h43c;
	10'd422 : sinewave = 12'h431;
	10'd423 : sinewave = 12'h427;
	10'd424 : sinewave = 12'h41c;
	10'd425 : sinewave = 12'h411;
	10'd426 : sinewave = 12'h406;
	10'd427 : sinewave = 12'h3fb;
	10'd428 : sinewave = 12'h3f0;
	10'd429 : sinewave = 12'h3e6;
	10'd430 : sinewave = 12'h3db;
	10'd431 : sinewave = 12'h3d0;
	10'd432 : sinewave = 12'h3c4;
	10'd433 : sinewave = 12'h3b9;
	10'd434 : sinewave = 12'h3ae;
	10'd435 : sinewave = 12'h3a3;
	10'd436 : sinewave = 12'h398;
	10'd437 : sinewave = 12'h38d;
	10'd438 : sinewave = 12'h381;
	10'd439 : sinewave = 12'h376;
	10'd440 : sinewave = 12'h36b;
	10'd441 : sinewave = 12'h35f;
	10'd442 : sinewave = 12'h354;
	10'd443 : sinewave = 12'h348;
	10'd444 : sinewave = 12'h33d;
	10'd445 : sinewave = 12'h332;
	10'd446 : sinewave = 12'h326;
	10'd447 : sinewave = 12'h31a;
	10'd448 : sinewave = 12'h30f;
	10'd449 : sinewave = 12'h303;
	10'd450 : sinewave = 12'h2f8;
	10'd451 : sinewave = 12'h2ec;
	10'd452 : sinewave = 12'h2e0;
	10'd453 : sinewave = 12'h2d4;
	10'd454 : sinewave = 12'h2c9;
	10'd455 : sinewave = 12'h2bd;
	10'd456 : sinewave = 12'h2b1;
	10'd457 : sinewave = 12'h2a5;
	10'd458 : sinewave = 12'h299;
	10'd459 : sinewave = 12'h28e;
	10'd460 : sinewave = 12'h282;
	10'd461 : sinewave = 12'h276;
	10'd462 : sinewave = 12'h26a;
	10'd463 : sinewave = 12'h25e;
	10'd464 : sinewave = 12'h252;
	10'd465 : sinewave = 12'h246;
	10'd466 : sinewave = 12'h23a;
	10'd467 : sinewave = 12'h22e;
	10'd468 : sinewave = 12'h221;
	10'd469 : sinewave = 12'h215;
	10'd470 : sinewave = 12'h209;
	10'd471 : sinewave = 12'h1fd;
	10'd472 : sinewave = 12'h1f1;
	10'd473 : sinewave = 12'h1e5;
	10'd474 : sinewave = 12'h1d8;
	10'd475 : sinewave = 12'h1cc;
	10'd476 : sinewave = 12'h1c0;
	10'd477 : sinewave = 12'h1b4;
	10'd478 : sinewave = 12'h1a7;
	10'd479 : sinewave = 12'h19b;
	10'd480 : sinewave = 12'h18f;
	10'd481 : sinewave = 12'h183;
	10'd482 : sinewave = 12'h176;
	10'd483 : sinewave = 12'h16a;
	10'd484 : sinewave = 12'h15d;
	10'd485 : sinewave = 12'h151;
	10'd486 : sinewave = 12'h145;
	10'd487 : sinewave = 12'h138;
	10'd488 : sinewave = 12'h12c;
	10'd489 : sinewave = 12'h11f;
	10'd490 : sinewave = 12'h113;
	10'd491 : sinewave = 12'h107;
	10'd492 : sinewave = 12'hfa;
	10'd493 : sinewave = 12'hee;
	10'd494 : sinewave = 12'he1;
	10'd495 : sinewave = 12'hd5;
	10'd496 : sinewave = 12'hc8;
	10'd497 : sinewave = 12'hbc;
	10'd498 : sinewave = 12'haf;
	10'd499 : sinewave = 12'ha3;
	10'd500 : sinewave = 12'h96;
	10'd501 : sinewave = 12'h8a;
	10'd502 : sinewave = 12'h7d;
	10'd503 : sinewave = 12'h70;
	10'd504 : sinewave = 12'h64;
	10'd505 : sinewave = 12'h57;
	10'd506 : sinewave = 12'h4b;
	10'd507 : sinewave = 12'h3e;
	10'd508 : sinewave = 12'h32;
	10'd509 : sinewave = 12'h25;
	10'd510 : sinewave = 12'h19;
	10'd511 : sinewave = 12'h0c;
	10'd512 : sinewave = 12'h00;
	10'd513 : sinewave = 12'hff4;
	10'd514 : sinewave = 12'hfe7;
	10'd515 : sinewave = 12'hfdb;
	10'd516 : sinewave = 12'hfce;
	10'd517 : sinewave = 12'hfc2;
	10'd518 : sinewave = 12'hfb5;
	10'd519 : sinewave = 12'hfa9;
	10'd520 : sinewave = 12'hf9c;
	10'd521 : sinewave = 12'hf90;
	10'd522 : sinewave = 12'hf83;
	10'd523 : sinewave = 12'hf76;
	10'd524 : sinewave = 12'hf6a;
	10'd525 : sinewave = 12'hf5d;
	10'd526 : sinewave = 12'hf51;
	10'd527 : sinewave = 12'hf44;
	10'd528 : sinewave = 12'hf38;
	10'd529 : sinewave = 12'hf2b;
	10'd530 : sinewave = 12'hf1f;
	10'd531 : sinewave = 12'hf12;
	10'd532 : sinewave = 12'hf06;
	10'd533 : sinewave = 12'hef9;
	10'd534 : sinewave = 12'heed;
	10'd535 : sinewave = 12'hee1;
	10'd536 : sinewave = 12'hed4;
	10'd537 : sinewave = 12'hec8;
	10'd538 : sinewave = 12'hebb;
	10'd539 : sinewave = 12'heaf;
	10'd540 : sinewave = 12'hea3;
	10'd541 : sinewave = 12'he96;
	10'd542 : sinewave = 12'he8a;
	10'd543 : sinewave = 12'he7d;
	10'd544 : sinewave = 12'he71;
	10'd545 : sinewave = 12'he65;
	10'd546 : sinewave = 12'he59;
	10'd547 : sinewave = 12'he4c;
	10'd548 : sinewave = 12'he40;
	10'd549 : sinewave = 12'he34;
	10'd550 : sinewave = 12'he28;
	10'd551 : sinewave = 12'he1b;
	10'd552 : sinewave = 12'he0f;
	10'd553 : sinewave = 12'he03;
	10'd554 : sinewave = 12'hdf7;
	10'd555 : sinewave = 12'hdeb;
	10'd556 : sinewave = 12'hddf;
	10'd557 : sinewave = 12'hdd2;
	10'd558 : sinewave = 12'hdc6;
	10'd559 : sinewave = 12'hdba;
	10'd560 : sinewave = 12'hdae;
	10'd561 : sinewave = 12'hda2;
	10'd562 : sinewave = 12'hd96;
	10'd563 : sinewave = 12'hd8a;
	10'd564 : sinewave = 12'hd7e;
	10'd565 : sinewave = 12'hd72;
	10'd566 : sinewave = 12'hd67;
	10'd567 : sinewave = 12'hd5b;
	10'd568 : sinewave = 12'hd4f;
	10'd569 : sinewave = 12'hd43;
	10'd570 : sinewave = 12'hd37;
	10'd571 : sinewave = 12'hd2c;
	10'd572 : sinewave = 12'hd20;
	10'd573 : sinewave = 12'hd14;
	10'd574 : sinewave = 12'hd08;
	10'd575 : sinewave = 12'hcfd;
	10'd576 : sinewave = 12'hcf1;
	10'd577 : sinewave = 12'hce6;
	10'd578 : sinewave = 12'hcda;
	10'd579 : sinewave = 12'hcce;
	10'd580 : sinewave = 12'hcc3;
	10'd581 : sinewave = 12'hcb8;
	10'd582 : sinewave = 12'hcac;
	10'd583 : sinewave = 12'hca1;
	10'd584 : sinewave = 12'hc95;
	10'd585 : sinewave = 12'hc8a;
	10'd586 : sinewave = 12'hc7f;
	10'd587 : sinewave = 12'hc73;
	10'd588 : sinewave = 12'hc68;
	10'd589 : sinewave = 12'hc5d;
	10'd590 : sinewave = 12'hc52;
	10'd591 : sinewave = 12'hc47;
	10'd592 : sinewave = 12'hc3c;
	10'd593 : sinewave = 12'hc30;
	10'd594 : sinewave = 12'hc25;
	10'd595 : sinewave = 12'hc1a;
	10'd596 : sinewave = 12'hc10;
	10'd597 : sinewave = 12'hc05;
	10'd598 : sinewave = 12'hbfa;
	10'd599 : sinewave = 12'hbef;
	10'd600 : sinewave = 12'hbe4;
	10'd601 : sinewave = 12'hbd9;
	10'd602 : sinewave = 12'hbcf;
	10'd603 : sinewave = 12'hbc4;
	10'd604 : sinewave = 12'hbb9;
	10'd605 : sinewave = 12'hbaf;
	10'd606 : sinewave = 12'hba4;
	10'd607 : sinewave = 12'hb9a;
	10'd608 : sinewave = 12'hb8f;
	10'd609 : sinewave = 12'hb85;
	10'd610 : sinewave = 12'hb7a;
	10'd611 : sinewave = 12'hb70;
	10'd612 : sinewave = 12'hb66;
	10'd613 : sinewave = 12'hb5c;
	10'd614 : sinewave = 12'hb51;
	10'd615 : sinewave = 12'hb47;
	10'd616 : sinewave = 12'hb3d;
	10'd617 : sinewave = 12'hb33;
	10'd618 : sinewave = 12'hb29;
	10'd619 : sinewave = 12'hb1f;
	10'd620 : sinewave = 12'hb15;
	10'd621 : sinewave = 12'hb0b;
	10'd622 : sinewave = 12'hb01;
	10'd623 : sinewave = 12'haf8;
	10'd624 : sinewave = 12'haee;
	10'd625 : sinewave = 12'hae4;
	10'd626 : sinewave = 12'hadb;
	10'd627 : sinewave = 12'had1;
	10'd628 : sinewave = 12'hac7;
	10'd629 : sinewave = 12'habe;
	10'd630 : sinewave = 12'hab5;
	10'd631 : sinewave = 12'haab;
	10'd632 : sinewave = 12'haa2;
	10'd633 : sinewave = 12'ha99;
	10'd634 : sinewave = 12'ha8f;
	10'd635 : sinewave = 12'ha86;
	10'd636 : sinewave = 12'ha7d;
	10'd637 : sinewave = 12'ha74;
	10'd638 : sinewave = 12'ha6b;
	10'd639 : sinewave = 12'ha62;
	10'd640 : sinewave = 12'ha59;
	10'd641 : sinewave = 12'ha50;
	10'd642 : sinewave = 12'ha47;
	10'd643 : sinewave = 12'ha3f;
	10'd644 : sinewave = 12'ha36;
	10'd645 : sinewave = 12'ha2d;
	10'd646 : sinewave = 12'ha25;
	10'd647 : sinewave = 12'ha1c;
	10'd648 : sinewave = 12'ha14;
	10'd649 : sinewave = 12'ha0b;
	10'd650 : sinewave = 12'ha03;
	10'd651 : sinewave = 12'h9fb;
	10'd652 : sinewave = 12'h9f2;
	10'd653 : sinewave = 12'h9ea;
	10'd654 : sinewave = 12'h9e2;
	10'd655 : sinewave = 12'h9da;
	10'd656 : sinewave = 12'h9d2;
	10'd657 : sinewave = 12'h9ca;
	10'd658 : sinewave = 12'h9c2;
	10'd659 : sinewave = 12'h9bb;
	10'd660 : sinewave = 12'h9b3;
	10'd661 : sinewave = 12'h9ab;
	10'd662 : sinewave = 12'h9a3;
	10'd663 : sinewave = 12'h99c;
	10'd664 : sinewave = 12'h994;
	10'd665 : sinewave = 12'h98d;
	10'd666 : sinewave = 12'h985;
	10'd667 : sinewave = 12'h97e;
	10'd668 : sinewave = 12'h977;
	10'd669 : sinewave = 12'h970;
	10'd670 : sinewave = 12'h969;
	10'd671 : sinewave = 12'h961;
	10'd672 : sinewave = 12'h95a;
	10'd673 : sinewave = 12'h954;
	10'd674 : sinewave = 12'h94d;
	10'd675 : sinewave = 12'h946;
	10'd676 : sinewave = 12'h93f;
	10'd677 : sinewave = 12'h938;
	10'd678 : sinewave = 12'h932;
	10'd679 : sinewave = 12'h92b;
	10'd680 : sinewave = 12'h925;
	10'd681 : sinewave = 12'h91e;
	10'd682 : sinewave = 12'h918;
	10'd683 : sinewave = 12'h912;
	10'd684 : sinewave = 12'h90b;
	10'd685 : sinewave = 12'h905;
	10'd686 : sinewave = 12'h8ff;
	10'd687 : sinewave = 12'h8f9;
	10'd688 : sinewave = 12'h8f3;
	10'd689 : sinewave = 12'h8ed;
	10'd690 : sinewave = 12'h8e8;
	10'd691 : sinewave = 12'h8e2;
	10'd692 : sinewave = 12'h8dc;
	10'd693 : sinewave = 12'h8d6;
	10'd694 : sinewave = 12'h8d1;
	10'd695 : sinewave = 12'h8cb;
	10'd696 : sinewave = 12'h8c6;
	10'd697 : sinewave = 12'h8c1;
	10'd698 : sinewave = 12'h8bb;
	10'd699 : sinewave = 12'h8b6;
	10'd700 : sinewave = 12'h8b1;
	10'd701 : sinewave = 12'h8ac;
	10'd702 : sinewave = 12'h8a7;
	10'd703 : sinewave = 12'h8a2;
	10'd704 : sinewave = 12'h89d;
	10'd705 : sinewave = 12'h899;
	10'd706 : sinewave = 12'h894;
	10'd707 : sinewave = 12'h88f;
	10'd708 : sinewave = 12'h88b;
	10'd709 : sinewave = 12'h886;
	10'd710 : sinewave = 12'h882;
	10'd711 : sinewave = 12'h87d;
	10'd712 : sinewave = 12'h879;
	10'd713 : sinewave = 12'h875;
	10'd714 : sinewave = 12'h871;
	10'd715 : sinewave = 12'h86d;
	10'd716 : sinewave = 12'h869;
	10'd717 : sinewave = 12'h865;
	10'd718 : sinewave = 12'h861;
	10'd719 : sinewave = 12'h85d;
	10'd720 : sinewave = 12'h85a;
	10'd721 : sinewave = 12'h856;
	10'd722 : sinewave = 12'h852;
	10'd723 : sinewave = 12'h84f;
	10'd724 : sinewave = 12'h84c;
	10'd725 : sinewave = 12'h848;
	10'd726 : sinewave = 12'h845;
	10'd727 : sinewave = 12'h842;
	10'd728 : sinewave = 12'h83f;
	10'd729 : sinewave = 12'h83c;
	10'd730 : sinewave = 12'h839;
	10'd731 : sinewave = 12'h836;
	10'd732 : sinewave = 12'h833;
	10'd733 : sinewave = 12'h831;
	10'd734 : sinewave = 12'h82e;
	10'd735 : sinewave = 12'h82b;
	10'd736 : sinewave = 12'h829;
	10'd737 : sinewave = 12'h826;
	10'd738 : sinewave = 12'h824;
	10'd739 : sinewave = 12'h822;
	10'd740 : sinewave = 12'h820;
	10'd741 : sinewave = 12'h81e;
	10'd742 : sinewave = 12'h81b;
	10'd743 : sinewave = 12'h81a;
	10'd744 : sinewave = 12'h818;
	10'd745 : sinewave = 12'h816;
	10'd746 : sinewave = 12'h814;
	10'd747 : sinewave = 12'h812;
	10'd748 : sinewave = 12'h811;
	10'd749 : sinewave = 12'h80f;
	10'd750 : sinewave = 12'h80e;
	10'd751 : sinewave = 12'h80d;
	10'd752 : sinewave = 12'h80b;
	10'd753 : sinewave = 12'h80a;
	10'd754 : sinewave = 12'h809;
	10'd755 : sinewave = 12'h808;
	10'd756 : sinewave = 12'h807;
	10'd757 : sinewave = 12'h806;
	10'd758 : sinewave = 12'h805;
	10'd759 : sinewave = 12'h805;
	10'd760 : sinewave = 12'h804;
	10'd761 : sinewave = 12'h803;
	10'd762 : sinewave = 12'h803;
	10'd763 : sinewave = 12'h802;
	10'd764 : sinewave = 12'h802;
	10'd765 : sinewave = 12'h802;
	10'd766 : sinewave = 12'h802;
	10'd767 : sinewave = 12'h802;
	10'd768 : sinewave = 12'h801;
	10'd769 : sinewave = 12'h802;
	10'd770 : sinewave = 12'h802;
	10'd771 : sinewave = 12'h802;
	10'd772 : sinewave = 12'h802;
	10'd773 : sinewave = 12'h802;
	10'd774 : sinewave = 12'h803;
	10'd775 : sinewave = 12'h803;
	10'd776 : sinewave = 12'h804;
	10'd777 : sinewave = 12'h805;
	10'd778 : sinewave = 12'h805;
	10'd779 : sinewave = 12'h806;
	10'd780 : sinewave = 12'h807;
	10'd781 : sinewave = 12'h808;
	10'd782 : sinewave = 12'h809;
	10'd783 : sinewave = 12'h80a;
	10'd784 : sinewave = 12'h80b;
	10'd785 : sinewave = 12'h80d;
	10'd786 : sinewave = 12'h80e;
	10'd787 : sinewave = 12'h80f;
	10'd788 : sinewave = 12'h811;
	10'd789 : sinewave = 12'h812;
	10'd790 : sinewave = 12'h814;
	10'd791 : sinewave = 12'h816;
	10'd792 : sinewave = 12'h818;
	10'd793 : sinewave = 12'h81a;
	10'd794 : sinewave = 12'h81b;
	10'd795 : sinewave = 12'h81e;
	10'd796 : sinewave = 12'h820;
	10'd797 : sinewave = 12'h822;
	10'd798 : sinewave = 12'h824;
	10'd799 : sinewave = 12'h826;
	10'd800 : sinewave = 12'h829;
	10'd801 : sinewave = 12'h82b;
	10'd802 : sinewave = 12'h82e;
	10'd803 : sinewave = 12'h831;
	10'd804 : sinewave = 12'h833;
	10'd805 : sinewave = 12'h836;
	10'd806 : sinewave = 12'h839;
	10'd807 : sinewave = 12'h83c;
	10'd808 : sinewave = 12'h83f;
	10'd809 : sinewave = 12'h842;
	10'd810 : sinewave = 12'h845;
	10'd811 : sinewave = 12'h848;
	10'd812 : sinewave = 12'h84c;
	10'd813 : sinewave = 12'h84f;
	10'd814 : sinewave = 12'h852;
	10'd815 : sinewave = 12'h856;
	10'd816 : sinewave = 12'h85a;
	10'd817 : sinewave = 12'h85d;
	10'd818 : sinewave = 12'h861;
	10'd819 : sinewave = 12'h865;
	10'd820 : sinewave = 12'h869;
	10'd821 : sinewave = 12'h86d;
	10'd822 : sinewave = 12'h871;
	10'd823 : sinewave = 12'h875;
	10'd824 : sinewave = 12'h879;
	10'd825 : sinewave = 12'h87d;
	10'd826 : sinewave = 12'h882;
	10'd827 : sinewave = 12'h886;
	10'd828 : sinewave = 12'h88b;
	10'd829 : sinewave = 12'h88f;
	10'd830 : sinewave = 12'h894;
	10'd831 : sinewave = 12'h899;
	10'd832 : sinewave = 12'h89d;
	10'd833 : sinewave = 12'h8a2;
	10'd834 : sinewave = 12'h8a7;
	10'd835 : sinewave = 12'h8ac;
	10'd836 : sinewave = 12'h8b1;
	10'd837 : sinewave = 12'h8b6;
	10'd838 : sinewave = 12'h8bb;
	10'd839 : sinewave = 12'h8c1;
	10'd840 : sinewave = 12'h8c6;
	10'd841 : sinewave = 12'h8cb;
	10'd842 : sinewave = 12'h8d1;
	10'd843 : sinewave = 12'h8d6;
	10'd844 : sinewave = 12'h8dc;
	10'd845 : sinewave = 12'h8e2;
	10'd846 : sinewave = 12'h8e8;
	10'd847 : sinewave = 12'h8ed;
	10'd848 : sinewave = 12'h8f3;
	10'd849 : sinewave = 12'h8f9;
	10'd850 : sinewave = 12'h8ff;
	10'd851 : sinewave = 12'h905;
	10'd852 : sinewave = 12'h90b;
	10'd853 : sinewave = 12'h912;
	10'd854 : sinewave = 12'h918;
	10'd855 : sinewave = 12'h91e;
	10'd856 : sinewave = 12'h925;
	10'd857 : sinewave = 12'h92b;
	10'd858 : sinewave = 12'h932;
	10'd859 : sinewave = 12'h938;
	10'd860 : sinewave = 12'h93f;
	10'd861 : sinewave = 12'h946;
	10'd862 : sinewave = 12'h94d;
	10'd863 : sinewave = 12'h954;
	10'd864 : sinewave = 12'h95a;
	10'd865 : sinewave = 12'h961;
	10'd866 : sinewave = 12'h969;
	10'd867 : sinewave = 12'h970;
	10'd868 : sinewave = 12'h977;
	10'd869 : sinewave = 12'h97e;
	10'd870 : sinewave = 12'h985;
	10'd871 : sinewave = 12'h98d;
	10'd872 : sinewave = 12'h994;
	10'd873 : sinewave = 12'h99c;
	10'd874 : sinewave = 12'h9a3;
	10'd875 : sinewave = 12'h9ab;
	10'd876 : sinewave = 12'h9b3;
	10'd877 : sinewave = 12'h9bb;
	10'd878 : sinewave = 12'h9c2;
	10'd879 : sinewave = 12'h9ca;
	10'd880 : sinewave = 12'h9d2;
	10'd881 : sinewave = 12'h9da;
	10'd882 : sinewave = 12'h9e2;
	10'd883 : sinewave = 12'h9ea;
	10'd884 : sinewave = 12'h9f2;
	10'd885 : sinewave = 12'h9fb;
	10'd886 : sinewave = 12'ha03;
	10'd887 : sinewave = 12'ha0b;
	10'd888 : sinewave = 12'ha14;
	10'd889 : sinewave = 12'ha1c;
	10'd890 : sinewave = 12'ha25;
	10'd891 : sinewave = 12'ha2d;
	10'd892 : sinewave = 12'ha36;
	10'd893 : sinewave = 12'ha3f;
	10'd894 : sinewave = 12'ha47;
	10'd895 : sinewave = 12'ha50;
	10'd896 : sinewave = 12'ha59;
	10'd897 : sinewave = 12'ha62;
	10'd898 : sinewave = 12'ha6b;
	10'd899 : sinewave = 12'ha74;
	10'd900 : sinewave = 12'ha7d;
	10'd901 : sinewave = 12'ha86;
	10'd902 : sinewave = 12'ha8f;
	10'd903 : sinewave = 12'ha99;
	10'd904 : sinewave = 12'haa2;
	10'd905 : sinewave = 12'haab;
	10'd906 : sinewave = 12'hab5;
	10'd907 : sinewave = 12'habe;
	10'd908 : sinewave = 12'hac7;
	10'd909 : sinewave = 12'had1;
	10'd910 : sinewave = 12'hadb;
	10'd911 : sinewave = 12'hae4;
	10'd912 : sinewave = 12'haee;
	10'd913 : sinewave = 12'haf8;
	10'd914 : sinewave = 12'hb01;
	10'd915 : sinewave = 12'hb0b;
	10'd916 : sinewave = 12'hb15;
	10'd917 : sinewave = 12'hb1f;
	10'd918 : sinewave = 12'hb29;
	10'd919 : sinewave = 12'hb33;
	10'd920 : sinewave = 12'hb3d;
	10'd921 : sinewave = 12'hb47;
	10'd922 : sinewave = 12'hb51;
	10'd923 : sinewave = 12'hb5c;
	10'd924 : sinewave = 12'hb66;
	10'd925 : sinewave = 12'hb70;
	10'd926 : sinewave = 12'hb7a;
	10'd927 : sinewave = 12'hb85;
	10'd928 : sinewave = 12'hb8f;
	10'd929 : sinewave = 12'hb9a;
	10'd930 : sinewave = 12'hba4;
	10'd931 : sinewave = 12'hbaf;
	10'd932 : sinewave = 12'hbb9;
	10'd933 : sinewave = 12'hbc4;
	10'd934 : sinewave = 12'hbcf;
	10'd935 : sinewave = 12'hbd9;
	10'd936 : sinewave = 12'hbe4;
	10'd937 : sinewave = 12'hbef;
	10'd938 : sinewave = 12'hbfa;
	10'd939 : sinewave = 12'hc05;
	10'd940 : sinewave = 12'hc10;
	10'd941 : sinewave = 12'hc1a;
	10'd942 : sinewave = 12'hc25;
	10'd943 : sinewave = 12'hc30;
	10'd944 : sinewave = 12'hc3c;
	10'd945 : sinewave = 12'hc47;
	10'd946 : sinewave = 12'hc52;
	10'd947 : sinewave = 12'hc5d;
	10'd948 : sinewave = 12'hc68;
	10'd949 : sinewave = 12'hc73;
	10'd950 : sinewave = 12'hc7f;
	10'd951 : sinewave = 12'hc8a;
	10'd952 : sinewave = 12'hc95;
	10'd953 : sinewave = 12'hca1;
	10'd954 : sinewave = 12'hcac;
	10'd955 : sinewave = 12'hcb8;
	10'd956 : sinewave = 12'hcc3;
	10'd957 : sinewave = 12'hcce;
	10'd958 : sinewave = 12'hcda;
	10'd959 : sinewave = 12'hce6;
	10'd960 : sinewave = 12'hcf1;
	10'd961 : sinewave = 12'hcfd;
	10'd962 : sinewave = 12'hd08;
	10'd963 : sinewave = 12'hd14;
	10'd964 : sinewave = 12'hd20;
	10'd965 : sinewave = 12'hd2c;
	10'd966 : sinewave = 12'hd37;
	10'd967 : sinewave = 12'hd43;
	10'd968 : sinewave = 12'hd4f;
	10'd969 : sinewave = 12'hd5b;
	10'd970 : sinewave = 12'hd67;
	10'd971 : sinewave = 12'hd72;
	10'd972 : sinewave = 12'hd7e;
	10'd973 : sinewave = 12'hd8a;
	10'd974 : sinewave = 12'hd96;
	10'd975 : sinewave = 12'hda2;
	10'd976 : sinewave = 12'hdae;
	10'd977 : sinewave = 12'hdba;
	10'd978 : sinewave = 12'hdc6;
	10'd979 : sinewave = 12'hdd2;
	10'd980 : sinewave = 12'hddf;
	10'd981 : sinewave = 12'hdeb;
	10'd982 : sinewave = 12'hdf7;
	10'd983 : sinewave = 12'he03;
	10'd984 : sinewave = 12'he0f;
	10'd985 : sinewave = 12'he1b;
	10'd986 : sinewave = 12'he28;
	10'd987 : sinewave = 12'he34;
	10'd988 : sinewave = 12'he40;
	10'd989 : sinewave = 12'he4c;
	10'd990 : sinewave = 12'he59;
	10'd991 : sinewave = 12'he65;
	10'd992 : sinewave = 12'he71;
	10'd993 : sinewave = 12'he7d;
	10'd994 : sinewave = 12'he8a;
	10'd995 : sinewave = 12'he96;
	10'd996 : sinewave = 12'hea3;
	10'd997 : sinewave = 12'heaf;
	10'd998 : sinewave = 12'hebb;
	10'd999 : sinewave = 12'hec8;
	10'd1000: sinewave = 12'hed4;
	10'd1001: sinewave = 12'hee1;
	10'd1002: sinewave = 12'heed;
	10'd1003: sinewave = 12'hef9;
	10'd1004: sinewave = 12'hf06;
	10'd1005: sinewave = 12'hf12;
	10'd1006: sinewave = 12'hf1f;
	10'd1007: sinewave = 12'hf2b;
	10'd1008: sinewave = 12'hf38;
	10'd1009: sinewave = 12'hf44;
	10'd1010: sinewave = 12'hf51;
	10'd1011: sinewave = 12'hf5d;
	10'd1012: sinewave = 12'hf6a;
	10'd1013: sinewave = 12'hf76;
	10'd1014: sinewave = 12'hf83;
	10'd1015: sinewave = 12'hf90;
	10'd1016: sinewave = 12'hf9c;
	10'd1017: sinewave = 12'hfa9;
	10'd1018: sinewave = 12'hfb5;
	10'd1019: sinewave = 12'hfc2;
	10'd1020: sinewave = 12'hfce;
	10'd1021: sinewave = 12'hfdb;
	10'd1022: sinewave = 12'hfe7;
	10'd1023: sinewave = 12'hff4;
	endcase

end

endmodule
